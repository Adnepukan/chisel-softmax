module PipelineHsk(
  input   clock,
  input   reset,
  input   io_validPre,
  output  io_readyPre,
  input   io_lastPre,
  output  io_validNxt,
  input   io_readyNxt,
  output  io_regen_0,
  output  io_regen_1,
  output  io_lastNxt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  valid_1_r; // @[Reg.scala 28:20]
  reg  valid_2_r; // @[Reg.scala 28:20]
  wire  ready_1 = io_readyNxt | ~valid_2_r; // @[pipelinehsk.scala 24:32]
  wire  ready_0 = ready_1 | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  reg  last_1_r; // @[Reg.scala 28:20]
  reg  last_2_r; // @[Reg.scala 28:20]
  assign io_readyPre = ready_1 | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  assign io_validNxt = valid_2_r; // @[pipelinehsk.scala 17:21 22:20]
  assign io_regen_0 = io_validPre & ready_0; // @[pipelinehsk.scala 25:33]
  assign io_regen_1 = valid_1_r & ready_1; // @[pipelinehsk.scala 25:33]
  assign io_lastNxt = last_2_r; // @[pipelinehsk.scala 19:20 23:19]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_0) begin // @[Reg.scala 28:20]
      valid_1_r <= io_validPre;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_2_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_1) begin // @[Reg.scala 28:20]
      valid_2_r <= valid_1_r;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_0) begin // @[Reg.scala 28:20]
      last_1_r <= io_lastPre;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_2_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_1) begin // @[Reg.scala 28:20]
      last_2_r <= last_1_r;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_1_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_2_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  last_1_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  last_2_r = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid_1_r = 1'h0;
  end
  if (reset) begin
    valid_2_r = 1'h0;
  end
  if (reset) begin
    last_1_r = 1'h0;
  end
  if (reset) begin
    last_2_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Exponent(
  input        clock,
  input        reset,
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_x_0,
  input  [7:0] io_input_bits_x_1,
  input  [7:0] io_input_bits_x_2,
  input  [7:0] io_input_bits_x_3,
  input  [7:0] io_input_bits_x_4,
  input  [7:0] io_input_bits_x_5,
  input  [7:0] io_input_bits_x_6,
  input  [7:0] io_input_bits_x_7,
  input  [7:0] io_input_bits_x_8,
  input  [7:0] io_input_bits_x_9,
  input  [7:0] io_input_bits_x_10,
  input  [7:0] io_input_bits_x_11,
  input  [7:0] io_input_bits_x_12,
  input  [7:0] io_input_bits_x_13,
  input  [7:0] io_input_bits_x_14,
  input  [7:0] io_input_bits_x_15,
  input        io_input_bits_last,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_x_0,
  output [7:0] io_output_bits_x_1,
  output [7:0] io_output_bits_x_2,
  output [7:0] io_output_bits_x_3,
  output [7:0] io_output_bits_x_4,
  output [7:0] io_output_bits_x_5,
  output [7:0] io_output_bits_x_6,
  output [7:0] io_output_bits_x_7,
  output [7:0] io_output_bits_x_8,
  output [7:0] io_output_bits_x_9,
  output [7:0] io_output_bits_x_10,
  output [7:0] io_output_bits_x_11,
  output [7:0] io_output_bits_x_12,
  output [7:0] io_output_bits_x_13,
  output [7:0] io_output_bits_x_14,
  output [7:0] io_output_bits_x_15,
  output       io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  hsk_clock; // @[exponent.scala 20:21]
  wire  hsk_reset; // @[exponent.scala 20:21]
  wire  hsk_io_validPre; // @[exponent.scala 20:21]
  wire  hsk_io_readyPre; // @[exponent.scala 20:21]
  wire  hsk_io_lastPre; // @[exponent.scala 20:21]
  wire  hsk_io_validNxt; // @[exponent.scala 20:21]
  wire  hsk_io_readyNxt; // @[exponent.scala 20:21]
  wire  hsk_io_regen_0; // @[exponent.scala 20:21]
  wire  hsk_io_regen_1; // @[exponent.scala 20:21]
  wire  hsk_io_lastNxt; // @[exponent.scala 20:21]
  wire [12:0] _data1_T = $signed(io_input_bits_x_0) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_0; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_1 = $signed(io_input_bits_x_1) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_1; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_2 = $signed(io_input_bits_x_2) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_2; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_3 = $signed(io_input_bits_x_3) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_3; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_4 = $signed(io_input_bits_x_4) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_4; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_5 = $signed(io_input_bits_x_5) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_5; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_6 = $signed(io_input_bits_x_6) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_6; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_7 = $signed(io_input_bits_x_7) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_7; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_8 = $signed(io_input_bits_x_8) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_8; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_9 = $signed(io_input_bits_x_9) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_9; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_10 = $signed(io_input_bits_x_10) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_10; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_11 = $signed(io_input_bits_x_11) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_11; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_12 = $signed(io_input_bits_x_12) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_12; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_13 = $signed(io_input_bits_x_13) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_13; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_14 = $signed(io_input_bits_x_14) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_14; // @[Reg.scala 16:16]
  wire [12:0] _data1_T_15 = $signed(io_input_bits_x_15) * 5'shc; // @[exponent.scala 30:53]
  reg [12:0] data1_15; // @[Reg.scala 16:16]
  wire [5:0] data1Int_0 = data1_0[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_1 = data1_1[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_2 = data1_2[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_3 = data1_3[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_4 = data1_4[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_5 = data1_5[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_6 = data1_6[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_7 = data1_7[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_8 = data1_8[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_9 = data1_9[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_10 = data1_10[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_11 = data1_11[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_12 = data1_12[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_13 = data1_13[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_14 = data1_14[12:7]; // @[exponent.scala 31:31]
  wire [5:0] data1Int_15 = data1_15[12:7]; // @[exponent.scala 31:31]
  wire [6:0] data1Frac_0 = data1_0[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_1 = data1_1[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_2 = data1_2[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_3 = data1_3[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_4 = data1_4[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_5 = data1_5[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_6 = data1_6[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_7 = data1_7[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_8 = data1_8[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_9 = data1_9[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_10 = data1_10[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_11 = data1_11[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_12 = data1_12[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_13 = data1_13[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_14 = data1_14[6:0]; // @[exponent.scala 32:32]
  wire [6:0] data1Frac_15 = data1_15[6:0]; // @[exponent.scala 32:32]
  wire [7:0] _GEN_18 = 7'h2 == data1Frac_0 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_19 = 7'h3 == data1Frac_0 ? $signed(8'sh3f) : $signed(_GEN_18); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_20 = 7'h4 == data1Frac_0 ? $signed(8'sh3f) : $signed(_GEN_19); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_21 = 7'h5 == data1Frac_0 ? $signed(8'sh3e) : $signed(_GEN_20); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_22 = 7'h6 == data1Frac_0 ? $signed(8'sh3e) : $signed(_GEN_21); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_23 = 7'h7 == data1Frac_0 ? $signed(8'sh3e) : $signed(_GEN_22); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_24 = 7'h8 == data1Frac_0 ? $signed(8'sh3d) : $signed(_GEN_23); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_25 = 7'h9 == data1Frac_0 ? $signed(8'sh3d) : $signed(_GEN_24); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_26 = 7'ha == data1Frac_0 ? $signed(8'sh3d) : $signed(_GEN_25); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_27 = 7'hb == data1Frac_0 ? $signed(8'sh3c) : $signed(_GEN_26); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_28 = 7'hc == data1Frac_0 ? $signed(8'sh3c) : $signed(_GEN_27); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_29 = 7'hd == data1Frac_0 ? $signed(8'sh3c) : $signed(_GEN_28); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_30 = 7'he == data1Frac_0 ? $signed(8'sh3b) : $signed(_GEN_29); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_31 = 7'hf == data1Frac_0 ? $signed(8'sh3b) : $signed(_GEN_30); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_32 = 7'h10 == data1Frac_0 ? $signed(8'sh3b) : $signed(_GEN_31); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_33 = 7'h11 == data1Frac_0 ? $signed(8'sh3a) : $signed(_GEN_32); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_34 = 7'h12 == data1Frac_0 ? $signed(8'sh3a) : $signed(_GEN_33); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_35 = 7'h13 == data1Frac_0 ? $signed(8'sh3a) : $signed(_GEN_34); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_36 = 7'h14 == data1Frac_0 ? $signed(8'sh39) : $signed(_GEN_35); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_37 = 7'h15 == data1Frac_0 ? $signed(8'sh39) : $signed(_GEN_36); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_38 = 7'h16 == data1Frac_0 ? $signed(8'sh39) : $signed(_GEN_37); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_39 = 7'h17 == data1Frac_0 ? $signed(8'sh39) : $signed(_GEN_38); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_40 = 7'h18 == data1Frac_0 ? $signed(8'sh38) : $signed(_GEN_39); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_41 = 7'h19 == data1Frac_0 ? $signed(8'sh38) : $signed(_GEN_40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_42 = 7'h1a == data1Frac_0 ? $signed(8'sh38) : $signed(_GEN_41); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_43 = 7'h1b == data1Frac_0 ? $signed(8'sh37) : $signed(_GEN_42); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_44 = 7'h1c == data1Frac_0 ? $signed(8'sh37) : $signed(_GEN_43); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_45 = 7'h1d == data1Frac_0 ? $signed(8'sh37) : $signed(_GEN_44); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_46 = 7'h1e == data1Frac_0 ? $signed(8'sh36) : $signed(_GEN_45); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_47 = 7'h1f == data1Frac_0 ? $signed(8'sh36) : $signed(_GEN_46); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_48 = 7'h20 == data1Frac_0 ? $signed(8'sh36) : $signed(_GEN_47); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_49 = 7'h21 == data1Frac_0 ? $signed(8'sh36) : $signed(_GEN_48); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_50 = 7'h22 == data1Frac_0 ? $signed(8'sh35) : $signed(_GEN_49); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_51 = 7'h23 == data1Frac_0 ? $signed(8'sh35) : $signed(_GEN_50); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_52 = 7'h24 == data1Frac_0 ? $signed(8'sh35) : $signed(_GEN_51); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_53 = 7'h25 == data1Frac_0 ? $signed(8'sh34) : $signed(_GEN_52); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_54 = 7'h26 == data1Frac_0 ? $signed(8'sh34) : $signed(_GEN_53); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_55 = 7'h27 == data1Frac_0 ? $signed(8'sh34) : $signed(_GEN_54); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_56 = 7'h28 == data1Frac_0 ? $signed(8'sh34) : $signed(_GEN_55); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_57 = 7'h29 == data1Frac_0 ? $signed(8'sh33) : $signed(_GEN_56); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_58 = 7'h2a == data1Frac_0 ? $signed(8'sh33) : $signed(_GEN_57); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_59 = 7'h2b == data1Frac_0 ? $signed(8'sh33) : $signed(_GEN_58); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_60 = 7'h2c == data1Frac_0 ? $signed(8'sh32) : $signed(_GEN_59); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_61 = 7'h2d == data1Frac_0 ? $signed(8'sh32) : $signed(_GEN_60); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_62 = 7'h2e == data1Frac_0 ? $signed(8'sh32) : $signed(_GEN_61); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_63 = 7'h2f == data1Frac_0 ? $signed(8'sh32) : $signed(_GEN_62); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_64 = 7'h30 == data1Frac_0 ? $signed(8'sh31) : $signed(_GEN_63); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_65 = 7'h31 == data1Frac_0 ? $signed(8'sh31) : $signed(_GEN_64); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_66 = 7'h32 == data1Frac_0 ? $signed(8'sh31) : $signed(_GEN_65); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_67 = 7'h33 == data1Frac_0 ? $signed(8'sh31) : $signed(_GEN_66); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_68 = 7'h34 == data1Frac_0 ? $signed(8'sh30) : $signed(_GEN_67); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_69 = 7'h35 == data1Frac_0 ? $signed(8'sh30) : $signed(_GEN_68); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_70 = 7'h36 == data1Frac_0 ? $signed(8'sh30) : $signed(_GEN_69); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_71 = 7'h37 == data1Frac_0 ? $signed(8'sh30) : $signed(_GEN_70); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_72 = 7'h38 == data1Frac_0 ? $signed(8'sh2f) : $signed(_GEN_71); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_73 = 7'h39 == data1Frac_0 ? $signed(8'sh2f) : $signed(_GEN_72); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_74 = 7'h3a == data1Frac_0 ? $signed(8'sh2f) : $signed(_GEN_73); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_75 = 7'h3b == data1Frac_0 ? $signed(8'sh2e) : $signed(_GEN_74); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_76 = 7'h3c == data1Frac_0 ? $signed(8'sh2e) : $signed(_GEN_75); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_77 = 7'h3d == data1Frac_0 ? $signed(8'sh2e) : $signed(_GEN_76); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_78 = 7'h3e == data1Frac_0 ? $signed(8'sh2e) : $signed(_GEN_77); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_79 = 7'h3f == data1Frac_0 ? $signed(8'sh2e) : $signed(_GEN_78); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_80 = 7'h40 == data1Frac_0 ? $signed(8'sh2d) : $signed(_GEN_79); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_81 = 7'h41 == data1Frac_0 ? $signed(8'sh2d) : $signed(_GEN_80); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_82 = 7'h42 == data1Frac_0 ? $signed(8'sh2d) : $signed(_GEN_81); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_83 = 7'h43 == data1Frac_0 ? $signed(8'sh2d) : $signed(_GEN_82); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_84 = 7'h44 == data1Frac_0 ? $signed(8'sh2c) : $signed(_GEN_83); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_85 = 7'h45 == data1Frac_0 ? $signed(8'sh2c) : $signed(_GEN_84); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_86 = 7'h46 == data1Frac_0 ? $signed(8'sh2c) : $signed(_GEN_85); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_87 = 7'h47 == data1Frac_0 ? $signed(8'sh2c) : $signed(_GEN_86); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_88 = 7'h48 == data1Frac_0 ? $signed(8'sh2b) : $signed(_GEN_87); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_89 = 7'h49 == data1Frac_0 ? $signed(8'sh2b) : $signed(_GEN_88); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_90 = 7'h4a == data1Frac_0 ? $signed(8'sh2b) : $signed(_GEN_89); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_91 = 7'h4b == data1Frac_0 ? $signed(8'sh2b) : $signed(_GEN_90); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_92 = 7'h4c == data1Frac_0 ? $signed(8'sh2a) : $signed(_GEN_91); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_93 = 7'h4d == data1Frac_0 ? $signed(8'sh2a) : $signed(_GEN_92); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_94 = 7'h4e == data1Frac_0 ? $signed(8'sh2a) : $signed(_GEN_93); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_95 = 7'h4f == data1Frac_0 ? $signed(8'sh2a) : $signed(_GEN_94); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_96 = 7'h50 == data1Frac_0 ? $signed(8'sh29) : $signed(_GEN_95); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_97 = 7'h51 == data1Frac_0 ? $signed(8'sh29) : $signed(_GEN_96); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_98 = 7'h52 == data1Frac_0 ? $signed(8'sh29) : $signed(_GEN_97); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_99 = 7'h53 == data1Frac_0 ? $signed(8'sh29) : $signed(_GEN_98); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_100 = 7'h54 == data1Frac_0 ? $signed(8'sh29) : $signed(_GEN_99); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_101 = 7'h55 == data1Frac_0 ? $signed(8'sh28) : $signed(_GEN_100); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_102 = 7'h56 == data1Frac_0 ? $signed(8'sh28) : $signed(_GEN_101); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_103 = 7'h57 == data1Frac_0 ? $signed(8'sh28) : $signed(_GEN_102); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_104 = 7'h58 == data1Frac_0 ? $signed(8'sh28) : $signed(_GEN_103); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_105 = 7'h59 == data1Frac_0 ? $signed(8'sh28) : $signed(_GEN_104); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_106 = 7'h5a == data1Frac_0 ? $signed(8'sh27) : $signed(_GEN_105); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_107 = 7'h5b == data1Frac_0 ? $signed(8'sh27) : $signed(_GEN_106); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_108 = 7'h5c == data1Frac_0 ? $signed(8'sh27) : $signed(_GEN_107); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_109 = 7'h5d == data1Frac_0 ? $signed(8'sh27) : $signed(_GEN_108); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_110 = 7'h5e == data1Frac_0 ? $signed(8'sh26) : $signed(_GEN_109); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_111 = 7'h5f == data1Frac_0 ? $signed(8'sh26) : $signed(_GEN_110); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_112 = 7'h60 == data1Frac_0 ? $signed(8'sh26) : $signed(_GEN_111); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_113 = 7'h61 == data1Frac_0 ? $signed(8'sh26) : $signed(_GEN_112); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_114 = 7'h62 == data1Frac_0 ? $signed(8'sh26) : $signed(_GEN_113); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_115 = 7'h63 == data1Frac_0 ? $signed(8'sh25) : $signed(_GEN_114); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_116 = 7'h64 == data1Frac_0 ? $signed(8'sh25) : $signed(_GEN_115); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_117 = 7'h65 == data1Frac_0 ? $signed(8'sh25) : $signed(_GEN_116); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_118 = 7'h66 == data1Frac_0 ? $signed(8'sh25) : $signed(_GEN_117); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_119 = 7'h67 == data1Frac_0 ? $signed(8'sh25) : $signed(_GEN_118); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_120 = 7'h68 == data1Frac_0 ? $signed(8'sh24) : $signed(_GEN_119); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_121 = 7'h69 == data1Frac_0 ? $signed(8'sh24) : $signed(_GEN_120); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_122 = 7'h6a == data1Frac_0 ? $signed(8'sh24) : $signed(_GEN_121); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_123 = 7'h6b == data1Frac_0 ? $signed(8'sh24) : $signed(_GEN_122); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_124 = 7'h6c == data1Frac_0 ? $signed(8'sh24) : $signed(_GEN_123); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_125 = 7'h6d == data1Frac_0 ? $signed(8'sh23) : $signed(_GEN_124); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_126 = 7'h6e == data1Frac_0 ? $signed(8'sh23) : $signed(_GEN_125); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_127 = 7'h6f == data1Frac_0 ? $signed(8'sh23) : $signed(_GEN_126); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_128 = 7'h70 == data1Frac_0 ? $signed(8'sh23) : $signed(_GEN_127); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_129 = 7'h71 == data1Frac_0 ? $signed(8'sh23) : $signed(_GEN_128); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_130 = 7'h72 == data1Frac_0 ? $signed(8'sh23) : $signed(_GEN_129); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_131 = 7'h73 == data1Frac_0 ? $signed(8'sh22) : $signed(_GEN_130); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_132 = 7'h74 == data1Frac_0 ? $signed(8'sh22) : $signed(_GEN_131); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_133 = 7'h75 == data1Frac_0 ? $signed(8'sh22) : $signed(_GEN_132); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_134 = 7'h76 == data1Frac_0 ? $signed(8'sh22) : $signed(_GEN_133); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_135 = 7'h77 == data1Frac_0 ? $signed(8'sh22) : $signed(_GEN_134); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_136 = 7'h78 == data1Frac_0 ? $signed(8'sh21) : $signed(_GEN_135); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_137 = 7'h79 == data1Frac_0 ? $signed(8'sh21) : $signed(_GEN_136); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_138 = 7'h7a == data1Frac_0 ? $signed(8'sh21) : $signed(_GEN_137); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_139 = 7'h7b == data1Frac_0 ? $signed(8'sh21) : $signed(_GEN_138); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_140 = 7'h7c == data1Frac_0 ? $signed(8'sh21) : $signed(_GEN_139); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_141 = 7'h7d == data1Frac_0 ? $signed(8'sh21) : $signed(_GEN_140); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_142 = 7'h7e == data1Frac_0 ? $signed(8'sh20) : $signed(_GEN_141); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_143 = 7'h7f == data1Frac_0 ? $signed(8'sh20) : $signed(_GEN_142); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_2 = $signed(_GEN_143) >>> data1Int_0; // @[exponent.scala 38:85]
  reg [7:0] data2_0; // @[Reg.scala 16:16]
  wire [7:0] _GEN_147 = 7'h2 == data1Frac_1 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_148 = 7'h3 == data1Frac_1 ? $signed(8'sh3f) : $signed(_GEN_147); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_149 = 7'h4 == data1Frac_1 ? $signed(8'sh3f) : $signed(_GEN_148); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_150 = 7'h5 == data1Frac_1 ? $signed(8'sh3e) : $signed(_GEN_149); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_151 = 7'h6 == data1Frac_1 ? $signed(8'sh3e) : $signed(_GEN_150); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_152 = 7'h7 == data1Frac_1 ? $signed(8'sh3e) : $signed(_GEN_151); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_153 = 7'h8 == data1Frac_1 ? $signed(8'sh3d) : $signed(_GEN_152); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_154 = 7'h9 == data1Frac_1 ? $signed(8'sh3d) : $signed(_GEN_153); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_155 = 7'ha == data1Frac_1 ? $signed(8'sh3d) : $signed(_GEN_154); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_156 = 7'hb == data1Frac_1 ? $signed(8'sh3c) : $signed(_GEN_155); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_157 = 7'hc == data1Frac_1 ? $signed(8'sh3c) : $signed(_GEN_156); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_158 = 7'hd == data1Frac_1 ? $signed(8'sh3c) : $signed(_GEN_157); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_159 = 7'he == data1Frac_1 ? $signed(8'sh3b) : $signed(_GEN_158); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_160 = 7'hf == data1Frac_1 ? $signed(8'sh3b) : $signed(_GEN_159); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_161 = 7'h10 == data1Frac_1 ? $signed(8'sh3b) : $signed(_GEN_160); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_162 = 7'h11 == data1Frac_1 ? $signed(8'sh3a) : $signed(_GEN_161); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_163 = 7'h12 == data1Frac_1 ? $signed(8'sh3a) : $signed(_GEN_162); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_164 = 7'h13 == data1Frac_1 ? $signed(8'sh3a) : $signed(_GEN_163); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_165 = 7'h14 == data1Frac_1 ? $signed(8'sh39) : $signed(_GEN_164); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_166 = 7'h15 == data1Frac_1 ? $signed(8'sh39) : $signed(_GEN_165); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_167 = 7'h16 == data1Frac_1 ? $signed(8'sh39) : $signed(_GEN_166); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_168 = 7'h17 == data1Frac_1 ? $signed(8'sh39) : $signed(_GEN_167); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_169 = 7'h18 == data1Frac_1 ? $signed(8'sh38) : $signed(_GEN_168); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_170 = 7'h19 == data1Frac_1 ? $signed(8'sh38) : $signed(_GEN_169); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_171 = 7'h1a == data1Frac_1 ? $signed(8'sh38) : $signed(_GEN_170); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_172 = 7'h1b == data1Frac_1 ? $signed(8'sh37) : $signed(_GEN_171); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_173 = 7'h1c == data1Frac_1 ? $signed(8'sh37) : $signed(_GEN_172); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_174 = 7'h1d == data1Frac_1 ? $signed(8'sh37) : $signed(_GEN_173); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_175 = 7'h1e == data1Frac_1 ? $signed(8'sh36) : $signed(_GEN_174); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_176 = 7'h1f == data1Frac_1 ? $signed(8'sh36) : $signed(_GEN_175); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_177 = 7'h20 == data1Frac_1 ? $signed(8'sh36) : $signed(_GEN_176); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_178 = 7'h21 == data1Frac_1 ? $signed(8'sh36) : $signed(_GEN_177); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_179 = 7'h22 == data1Frac_1 ? $signed(8'sh35) : $signed(_GEN_178); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_180 = 7'h23 == data1Frac_1 ? $signed(8'sh35) : $signed(_GEN_179); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_181 = 7'h24 == data1Frac_1 ? $signed(8'sh35) : $signed(_GEN_180); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_182 = 7'h25 == data1Frac_1 ? $signed(8'sh34) : $signed(_GEN_181); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_183 = 7'h26 == data1Frac_1 ? $signed(8'sh34) : $signed(_GEN_182); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_184 = 7'h27 == data1Frac_1 ? $signed(8'sh34) : $signed(_GEN_183); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_185 = 7'h28 == data1Frac_1 ? $signed(8'sh34) : $signed(_GEN_184); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_186 = 7'h29 == data1Frac_1 ? $signed(8'sh33) : $signed(_GEN_185); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_187 = 7'h2a == data1Frac_1 ? $signed(8'sh33) : $signed(_GEN_186); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_188 = 7'h2b == data1Frac_1 ? $signed(8'sh33) : $signed(_GEN_187); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_189 = 7'h2c == data1Frac_1 ? $signed(8'sh32) : $signed(_GEN_188); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_190 = 7'h2d == data1Frac_1 ? $signed(8'sh32) : $signed(_GEN_189); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_191 = 7'h2e == data1Frac_1 ? $signed(8'sh32) : $signed(_GEN_190); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_192 = 7'h2f == data1Frac_1 ? $signed(8'sh32) : $signed(_GEN_191); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_193 = 7'h30 == data1Frac_1 ? $signed(8'sh31) : $signed(_GEN_192); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_194 = 7'h31 == data1Frac_1 ? $signed(8'sh31) : $signed(_GEN_193); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_195 = 7'h32 == data1Frac_1 ? $signed(8'sh31) : $signed(_GEN_194); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_196 = 7'h33 == data1Frac_1 ? $signed(8'sh31) : $signed(_GEN_195); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_197 = 7'h34 == data1Frac_1 ? $signed(8'sh30) : $signed(_GEN_196); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_198 = 7'h35 == data1Frac_1 ? $signed(8'sh30) : $signed(_GEN_197); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_199 = 7'h36 == data1Frac_1 ? $signed(8'sh30) : $signed(_GEN_198); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_200 = 7'h37 == data1Frac_1 ? $signed(8'sh30) : $signed(_GEN_199); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_201 = 7'h38 == data1Frac_1 ? $signed(8'sh2f) : $signed(_GEN_200); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_202 = 7'h39 == data1Frac_1 ? $signed(8'sh2f) : $signed(_GEN_201); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_203 = 7'h3a == data1Frac_1 ? $signed(8'sh2f) : $signed(_GEN_202); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_204 = 7'h3b == data1Frac_1 ? $signed(8'sh2e) : $signed(_GEN_203); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_205 = 7'h3c == data1Frac_1 ? $signed(8'sh2e) : $signed(_GEN_204); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_206 = 7'h3d == data1Frac_1 ? $signed(8'sh2e) : $signed(_GEN_205); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_207 = 7'h3e == data1Frac_1 ? $signed(8'sh2e) : $signed(_GEN_206); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_208 = 7'h3f == data1Frac_1 ? $signed(8'sh2e) : $signed(_GEN_207); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_209 = 7'h40 == data1Frac_1 ? $signed(8'sh2d) : $signed(_GEN_208); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_210 = 7'h41 == data1Frac_1 ? $signed(8'sh2d) : $signed(_GEN_209); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_211 = 7'h42 == data1Frac_1 ? $signed(8'sh2d) : $signed(_GEN_210); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_212 = 7'h43 == data1Frac_1 ? $signed(8'sh2d) : $signed(_GEN_211); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_213 = 7'h44 == data1Frac_1 ? $signed(8'sh2c) : $signed(_GEN_212); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_214 = 7'h45 == data1Frac_1 ? $signed(8'sh2c) : $signed(_GEN_213); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_215 = 7'h46 == data1Frac_1 ? $signed(8'sh2c) : $signed(_GEN_214); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_216 = 7'h47 == data1Frac_1 ? $signed(8'sh2c) : $signed(_GEN_215); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_217 = 7'h48 == data1Frac_1 ? $signed(8'sh2b) : $signed(_GEN_216); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_218 = 7'h49 == data1Frac_1 ? $signed(8'sh2b) : $signed(_GEN_217); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_219 = 7'h4a == data1Frac_1 ? $signed(8'sh2b) : $signed(_GEN_218); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_220 = 7'h4b == data1Frac_1 ? $signed(8'sh2b) : $signed(_GEN_219); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_221 = 7'h4c == data1Frac_1 ? $signed(8'sh2a) : $signed(_GEN_220); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_222 = 7'h4d == data1Frac_1 ? $signed(8'sh2a) : $signed(_GEN_221); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_223 = 7'h4e == data1Frac_1 ? $signed(8'sh2a) : $signed(_GEN_222); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_224 = 7'h4f == data1Frac_1 ? $signed(8'sh2a) : $signed(_GEN_223); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_225 = 7'h50 == data1Frac_1 ? $signed(8'sh29) : $signed(_GEN_224); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_226 = 7'h51 == data1Frac_1 ? $signed(8'sh29) : $signed(_GEN_225); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_227 = 7'h52 == data1Frac_1 ? $signed(8'sh29) : $signed(_GEN_226); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_228 = 7'h53 == data1Frac_1 ? $signed(8'sh29) : $signed(_GEN_227); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_229 = 7'h54 == data1Frac_1 ? $signed(8'sh29) : $signed(_GEN_228); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_230 = 7'h55 == data1Frac_1 ? $signed(8'sh28) : $signed(_GEN_229); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_231 = 7'h56 == data1Frac_1 ? $signed(8'sh28) : $signed(_GEN_230); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_232 = 7'h57 == data1Frac_1 ? $signed(8'sh28) : $signed(_GEN_231); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_233 = 7'h58 == data1Frac_1 ? $signed(8'sh28) : $signed(_GEN_232); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_234 = 7'h59 == data1Frac_1 ? $signed(8'sh28) : $signed(_GEN_233); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_235 = 7'h5a == data1Frac_1 ? $signed(8'sh27) : $signed(_GEN_234); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_236 = 7'h5b == data1Frac_1 ? $signed(8'sh27) : $signed(_GEN_235); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_237 = 7'h5c == data1Frac_1 ? $signed(8'sh27) : $signed(_GEN_236); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_238 = 7'h5d == data1Frac_1 ? $signed(8'sh27) : $signed(_GEN_237); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_239 = 7'h5e == data1Frac_1 ? $signed(8'sh26) : $signed(_GEN_238); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_240 = 7'h5f == data1Frac_1 ? $signed(8'sh26) : $signed(_GEN_239); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_241 = 7'h60 == data1Frac_1 ? $signed(8'sh26) : $signed(_GEN_240); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_242 = 7'h61 == data1Frac_1 ? $signed(8'sh26) : $signed(_GEN_241); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_243 = 7'h62 == data1Frac_1 ? $signed(8'sh26) : $signed(_GEN_242); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_244 = 7'h63 == data1Frac_1 ? $signed(8'sh25) : $signed(_GEN_243); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_245 = 7'h64 == data1Frac_1 ? $signed(8'sh25) : $signed(_GEN_244); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_246 = 7'h65 == data1Frac_1 ? $signed(8'sh25) : $signed(_GEN_245); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_247 = 7'h66 == data1Frac_1 ? $signed(8'sh25) : $signed(_GEN_246); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_248 = 7'h67 == data1Frac_1 ? $signed(8'sh25) : $signed(_GEN_247); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_249 = 7'h68 == data1Frac_1 ? $signed(8'sh24) : $signed(_GEN_248); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_250 = 7'h69 == data1Frac_1 ? $signed(8'sh24) : $signed(_GEN_249); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_251 = 7'h6a == data1Frac_1 ? $signed(8'sh24) : $signed(_GEN_250); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_252 = 7'h6b == data1Frac_1 ? $signed(8'sh24) : $signed(_GEN_251); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_253 = 7'h6c == data1Frac_1 ? $signed(8'sh24) : $signed(_GEN_252); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_254 = 7'h6d == data1Frac_1 ? $signed(8'sh23) : $signed(_GEN_253); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_255 = 7'h6e == data1Frac_1 ? $signed(8'sh23) : $signed(_GEN_254); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_256 = 7'h6f == data1Frac_1 ? $signed(8'sh23) : $signed(_GEN_255); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_257 = 7'h70 == data1Frac_1 ? $signed(8'sh23) : $signed(_GEN_256); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_258 = 7'h71 == data1Frac_1 ? $signed(8'sh23) : $signed(_GEN_257); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_259 = 7'h72 == data1Frac_1 ? $signed(8'sh23) : $signed(_GEN_258); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_260 = 7'h73 == data1Frac_1 ? $signed(8'sh22) : $signed(_GEN_259); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_261 = 7'h74 == data1Frac_1 ? $signed(8'sh22) : $signed(_GEN_260); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_262 = 7'h75 == data1Frac_1 ? $signed(8'sh22) : $signed(_GEN_261); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_263 = 7'h76 == data1Frac_1 ? $signed(8'sh22) : $signed(_GEN_262); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_264 = 7'h77 == data1Frac_1 ? $signed(8'sh22) : $signed(_GEN_263); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_265 = 7'h78 == data1Frac_1 ? $signed(8'sh21) : $signed(_GEN_264); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_266 = 7'h79 == data1Frac_1 ? $signed(8'sh21) : $signed(_GEN_265); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_267 = 7'h7a == data1Frac_1 ? $signed(8'sh21) : $signed(_GEN_266); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_268 = 7'h7b == data1Frac_1 ? $signed(8'sh21) : $signed(_GEN_267); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_269 = 7'h7c == data1Frac_1 ? $signed(8'sh21) : $signed(_GEN_268); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_270 = 7'h7d == data1Frac_1 ? $signed(8'sh21) : $signed(_GEN_269); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_271 = 7'h7e == data1Frac_1 ? $signed(8'sh20) : $signed(_GEN_270); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_272 = 7'h7f == data1Frac_1 ? $signed(8'sh20) : $signed(_GEN_271); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_5 = $signed(_GEN_272) >>> data1Int_1; // @[exponent.scala 38:85]
  reg [7:0] data2_1; // @[Reg.scala 16:16]
  wire [7:0] _GEN_276 = 7'h2 == data1Frac_2 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_277 = 7'h3 == data1Frac_2 ? $signed(8'sh3f) : $signed(_GEN_276); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_278 = 7'h4 == data1Frac_2 ? $signed(8'sh3f) : $signed(_GEN_277); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_279 = 7'h5 == data1Frac_2 ? $signed(8'sh3e) : $signed(_GEN_278); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_280 = 7'h6 == data1Frac_2 ? $signed(8'sh3e) : $signed(_GEN_279); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_281 = 7'h7 == data1Frac_2 ? $signed(8'sh3e) : $signed(_GEN_280); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_282 = 7'h8 == data1Frac_2 ? $signed(8'sh3d) : $signed(_GEN_281); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_283 = 7'h9 == data1Frac_2 ? $signed(8'sh3d) : $signed(_GEN_282); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_284 = 7'ha == data1Frac_2 ? $signed(8'sh3d) : $signed(_GEN_283); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_285 = 7'hb == data1Frac_2 ? $signed(8'sh3c) : $signed(_GEN_284); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_286 = 7'hc == data1Frac_2 ? $signed(8'sh3c) : $signed(_GEN_285); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_287 = 7'hd == data1Frac_2 ? $signed(8'sh3c) : $signed(_GEN_286); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_288 = 7'he == data1Frac_2 ? $signed(8'sh3b) : $signed(_GEN_287); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_289 = 7'hf == data1Frac_2 ? $signed(8'sh3b) : $signed(_GEN_288); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_290 = 7'h10 == data1Frac_2 ? $signed(8'sh3b) : $signed(_GEN_289); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_291 = 7'h11 == data1Frac_2 ? $signed(8'sh3a) : $signed(_GEN_290); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_292 = 7'h12 == data1Frac_2 ? $signed(8'sh3a) : $signed(_GEN_291); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_293 = 7'h13 == data1Frac_2 ? $signed(8'sh3a) : $signed(_GEN_292); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_294 = 7'h14 == data1Frac_2 ? $signed(8'sh39) : $signed(_GEN_293); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_295 = 7'h15 == data1Frac_2 ? $signed(8'sh39) : $signed(_GEN_294); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_296 = 7'h16 == data1Frac_2 ? $signed(8'sh39) : $signed(_GEN_295); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_297 = 7'h17 == data1Frac_2 ? $signed(8'sh39) : $signed(_GEN_296); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_298 = 7'h18 == data1Frac_2 ? $signed(8'sh38) : $signed(_GEN_297); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_299 = 7'h19 == data1Frac_2 ? $signed(8'sh38) : $signed(_GEN_298); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_300 = 7'h1a == data1Frac_2 ? $signed(8'sh38) : $signed(_GEN_299); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_301 = 7'h1b == data1Frac_2 ? $signed(8'sh37) : $signed(_GEN_300); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_302 = 7'h1c == data1Frac_2 ? $signed(8'sh37) : $signed(_GEN_301); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_303 = 7'h1d == data1Frac_2 ? $signed(8'sh37) : $signed(_GEN_302); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_304 = 7'h1e == data1Frac_2 ? $signed(8'sh36) : $signed(_GEN_303); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_305 = 7'h1f == data1Frac_2 ? $signed(8'sh36) : $signed(_GEN_304); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_306 = 7'h20 == data1Frac_2 ? $signed(8'sh36) : $signed(_GEN_305); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_307 = 7'h21 == data1Frac_2 ? $signed(8'sh36) : $signed(_GEN_306); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_308 = 7'h22 == data1Frac_2 ? $signed(8'sh35) : $signed(_GEN_307); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_309 = 7'h23 == data1Frac_2 ? $signed(8'sh35) : $signed(_GEN_308); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_310 = 7'h24 == data1Frac_2 ? $signed(8'sh35) : $signed(_GEN_309); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_311 = 7'h25 == data1Frac_2 ? $signed(8'sh34) : $signed(_GEN_310); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_312 = 7'h26 == data1Frac_2 ? $signed(8'sh34) : $signed(_GEN_311); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_313 = 7'h27 == data1Frac_2 ? $signed(8'sh34) : $signed(_GEN_312); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_314 = 7'h28 == data1Frac_2 ? $signed(8'sh34) : $signed(_GEN_313); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_315 = 7'h29 == data1Frac_2 ? $signed(8'sh33) : $signed(_GEN_314); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_316 = 7'h2a == data1Frac_2 ? $signed(8'sh33) : $signed(_GEN_315); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_317 = 7'h2b == data1Frac_2 ? $signed(8'sh33) : $signed(_GEN_316); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_318 = 7'h2c == data1Frac_2 ? $signed(8'sh32) : $signed(_GEN_317); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_319 = 7'h2d == data1Frac_2 ? $signed(8'sh32) : $signed(_GEN_318); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_320 = 7'h2e == data1Frac_2 ? $signed(8'sh32) : $signed(_GEN_319); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_321 = 7'h2f == data1Frac_2 ? $signed(8'sh32) : $signed(_GEN_320); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_322 = 7'h30 == data1Frac_2 ? $signed(8'sh31) : $signed(_GEN_321); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_323 = 7'h31 == data1Frac_2 ? $signed(8'sh31) : $signed(_GEN_322); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_324 = 7'h32 == data1Frac_2 ? $signed(8'sh31) : $signed(_GEN_323); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_325 = 7'h33 == data1Frac_2 ? $signed(8'sh31) : $signed(_GEN_324); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_326 = 7'h34 == data1Frac_2 ? $signed(8'sh30) : $signed(_GEN_325); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_327 = 7'h35 == data1Frac_2 ? $signed(8'sh30) : $signed(_GEN_326); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_328 = 7'h36 == data1Frac_2 ? $signed(8'sh30) : $signed(_GEN_327); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_329 = 7'h37 == data1Frac_2 ? $signed(8'sh30) : $signed(_GEN_328); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_330 = 7'h38 == data1Frac_2 ? $signed(8'sh2f) : $signed(_GEN_329); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_331 = 7'h39 == data1Frac_2 ? $signed(8'sh2f) : $signed(_GEN_330); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_332 = 7'h3a == data1Frac_2 ? $signed(8'sh2f) : $signed(_GEN_331); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_333 = 7'h3b == data1Frac_2 ? $signed(8'sh2e) : $signed(_GEN_332); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_334 = 7'h3c == data1Frac_2 ? $signed(8'sh2e) : $signed(_GEN_333); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_335 = 7'h3d == data1Frac_2 ? $signed(8'sh2e) : $signed(_GEN_334); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_336 = 7'h3e == data1Frac_2 ? $signed(8'sh2e) : $signed(_GEN_335); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_337 = 7'h3f == data1Frac_2 ? $signed(8'sh2e) : $signed(_GEN_336); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_338 = 7'h40 == data1Frac_2 ? $signed(8'sh2d) : $signed(_GEN_337); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_339 = 7'h41 == data1Frac_2 ? $signed(8'sh2d) : $signed(_GEN_338); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_340 = 7'h42 == data1Frac_2 ? $signed(8'sh2d) : $signed(_GEN_339); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_341 = 7'h43 == data1Frac_2 ? $signed(8'sh2d) : $signed(_GEN_340); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_342 = 7'h44 == data1Frac_2 ? $signed(8'sh2c) : $signed(_GEN_341); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_343 = 7'h45 == data1Frac_2 ? $signed(8'sh2c) : $signed(_GEN_342); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_344 = 7'h46 == data1Frac_2 ? $signed(8'sh2c) : $signed(_GEN_343); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_345 = 7'h47 == data1Frac_2 ? $signed(8'sh2c) : $signed(_GEN_344); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_346 = 7'h48 == data1Frac_2 ? $signed(8'sh2b) : $signed(_GEN_345); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_347 = 7'h49 == data1Frac_2 ? $signed(8'sh2b) : $signed(_GEN_346); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_348 = 7'h4a == data1Frac_2 ? $signed(8'sh2b) : $signed(_GEN_347); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_349 = 7'h4b == data1Frac_2 ? $signed(8'sh2b) : $signed(_GEN_348); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_350 = 7'h4c == data1Frac_2 ? $signed(8'sh2a) : $signed(_GEN_349); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_351 = 7'h4d == data1Frac_2 ? $signed(8'sh2a) : $signed(_GEN_350); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_352 = 7'h4e == data1Frac_2 ? $signed(8'sh2a) : $signed(_GEN_351); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_353 = 7'h4f == data1Frac_2 ? $signed(8'sh2a) : $signed(_GEN_352); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_354 = 7'h50 == data1Frac_2 ? $signed(8'sh29) : $signed(_GEN_353); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_355 = 7'h51 == data1Frac_2 ? $signed(8'sh29) : $signed(_GEN_354); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_356 = 7'h52 == data1Frac_2 ? $signed(8'sh29) : $signed(_GEN_355); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_357 = 7'h53 == data1Frac_2 ? $signed(8'sh29) : $signed(_GEN_356); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_358 = 7'h54 == data1Frac_2 ? $signed(8'sh29) : $signed(_GEN_357); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_359 = 7'h55 == data1Frac_2 ? $signed(8'sh28) : $signed(_GEN_358); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_360 = 7'h56 == data1Frac_2 ? $signed(8'sh28) : $signed(_GEN_359); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_361 = 7'h57 == data1Frac_2 ? $signed(8'sh28) : $signed(_GEN_360); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_362 = 7'h58 == data1Frac_2 ? $signed(8'sh28) : $signed(_GEN_361); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_363 = 7'h59 == data1Frac_2 ? $signed(8'sh28) : $signed(_GEN_362); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_364 = 7'h5a == data1Frac_2 ? $signed(8'sh27) : $signed(_GEN_363); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_365 = 7'h5b == data1Frac_2 ? $signed(8'sh27) : $signed(_GEN_364); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_366 = 7'h5c == data1Frac_2 ? $signed(8'sh27) : $signed(_GEN_365); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_367 = 7'h5d == data1Frac_2 ? $signed(8'sh27) : $signed(_GEN_366); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_368 = 7'h5e == data1Frac_2 ? $signed(8'sh26) : $signed(_GEN_367); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_369 = 7'h5f == data1Frac_2 ? $signed(8'sh26) : $signed(_GEN_368); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_370 = 7'h60 == data1Frac_2 ? $signed(8'sh26) : $signed(_GEN_369); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_371 = 7'h61 == data1Frac_2 ? $signed(8'sh26) : $signed(_GEN_370); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_372 = 7'h62 == data1Frac_2 ? $signed(8'sh26) : $signed(_GEN_371); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_373 = 7'h63 == data1Frac_2 ? $signed(8'sh25) : $signed(_GEN_372); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_374 = 7'h64 == data1Frac_2 ? $signed(8'sh25) : $signed(_GEN_373); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_375 = 7'h65 == data1Frac_2 ? $signed(8'sh25) : $signed(_GEN_374); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_376 = 7'h66 == data1Frac_2 ? $signed(8'sh25) : $signed(_GEN_375); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_377 = 7'h67 == data1Frac_2 ? $signed(8'sh25) : $signed(_GEN_376); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_378 = 7'h68 == data1Frac_2 ? $signed(8'sh24) : $signed(_GEN_377); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_379 = 7'h69 == data1Frac_2 ? $signed(8'sh24) : $signed(_GEN_378); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_380 = 7'h6a == data1Frac_2 ? $signed(8'sh24) : $signed(_GEN_379); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_381 = 7'h6b == data1Frac_2 ? $signed(8'sh24) : $signed(_GEN_380); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_382 = 7'h6c == data1Frac_2 ? $signed(8'sh24) : $signed(_GEN_381); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_383 = 7'h6d == data1Frac_2 ? $signed(8'sh23) : $signed(_GEN_382); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_384 = 7'h6e == data1Frac_2 ? $signed(8'sh23) : $signed(_GEN_383); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_385 = 7'h6f == data1Frac_2 ? $signed(8'sh23) : $signed(_GEN_384); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_386 = 7'h70 == data1Frac_2 ? $signed(8'sh23) : $signed(_GEN_385); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_387 = 7'h71 == data1Frac_2 ? $signed(8'sh23) : $signed(_GEN_386); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_388 = 7'h72 == data1Frac_2 ? $signed(8'sh23) : $signed(_GEN_387); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_389 = 7'h73 == data1Frac_2 ? $signed(8'sh22) : $signed(_GEN_388); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_390 = 7'h74 == data1Frac_2 ? $signed(8'sh22) : $signed(_GEN_389); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_391 = 7'h75 == data1Frac_2 ? $signed(8'sh22) : $signed(_GEN_390); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_392 = 7'h76 == data1Frac_2 ? $signed(8'sh22) : $signed(_GEN_391); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_393 = 7'h77 == data1Frac_2 ? $signed(8'sh22) : $signed(_GEN_392); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_394 = 7'h78 == data1Frac_2 ? $signed(8'sh21) : $signed(_GEN_393); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_395 = 7'h79 == data1Frac_2 ? $signed(8'sh21) : $signed(_GEN_394); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_396 = 7'h7a == data1Frac_2 ? $signed(8'sh21) : $signed(_GEN_395); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_397 = 7'h7b == data1Frac_2 ? $signed(8'sh21) : $signed(_GEN_396); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_398 = 7'h7c == data1Frac_2 ? $signed(8'sh21) : $signed(_GEN_397); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_399 = 7'h7d == data1Frac_2 ? $signed(8'sh21) : $signed(_GEN_398); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_400 = 7'h7e == data1Frac_2 ? $signed(8'sh20) : $signed(_GEN_399); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_401 = 7'h7f == data1Frac_2 ? $signed(8'sh20) : $signed(_GEN_400); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_8 = $signed(_GEN_401) >>> data1Int_2; // @[exponent.scala 38:85]
  reg [7:0] data2_2; // @[Reg.scala 16:16]
  wire [7:0] _GEN_405 = 7'h2 == data1Frac_3 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_406 = 7'h3 == data1Frac_3 ? $signed(8'sh3f) : $signed(_GEN_405); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_407 = 7'h4 == data1Frac_3 ? $signed(8'sh3f) : $signed(_GEN_406); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_408 = 7'h5 == data1Frac_3 ? $signed(8'sh3e) : $signed(_GEN_407); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_409 = 7'h6 == data1Frac_3 ? $signed(8'sh3e) : $signed(_GEN_408); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_410 = 7'h7 == data1Frac_3 ? $signed(8'sh3e) : $signed(_GEN_409); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_411 = 7'h8 == data1Frac_3 ? $signed(8'sh3d) : $signed(_GEN_410); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_412 = 7'h9 == data1Frac_3 ? $signed(8'sh3d) : $signed(_GEN_411); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_413 = 7'ha == data1Frac_3 ? $signed(8'sh3d) : $signed(_GEN_412); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_414 = 7'hb == data1Frac_3 ? $signed(8'sh3c) : $signed(_GEN_413); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_415 = 7'hc == data1Frac_3 ? $signed(8'sh3c) : $signed(_GEN_414); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_416 = 7'hd == data1Frac_3 ? $signed(8'sh3c) : $signed(_GEN_415); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_417 = 7'he == data1Frac_3 ? $signed(8'sh3b) : $signed(_GEN_416); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_418 = 7'hf == data1Frac_3 ? $signed(8'sh3b) : $signed(_GEN_417); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_419 = 7'h10 == data1Frac_3 ? $signed(8'sh3b) : $signed(_GEN_418); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_420 = 7'h11 == data1Frac_3 ? $signed(8'sh3a) : $signed(_GEN_419); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_421 = 7'h12 == data1Frac_3 ? $signed(8'sh3a) : $signed(_GEN_420); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_422 = 7'h13 == data1Frac_3 ? $signed(8'sh3a) : $signed(_GEN_421); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_423 = 7'h14 == data1Frac_3 ? $signed(8'sh39) : $signed(_GEN_422); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_424 = 7'h15 == data1Frac_3 ? $signed(8'sh39) : $signed(_GEN_423); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_425 = 7'h16 == data1Frac_3 ? $signed(8'sh39) : $signed(_GEN_424); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_426 = 7'h17 == data1Frac_3 ? $signed(8'sh39) : $signed(_GEN_425); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_427 = 7'h18 == data1Frac_3 ? $signed(8'sh38) : $signed(_GEN_426); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_428 = 7'h19 == data1Frac_3 ? $signed(8'sh38) : $signed(_GEN_427); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_429 = 7'h1a == data1Frac_3 ? $signed(8'sh38) : $signed(_GEN_428); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_430 = 7'h1b == data1Frac_3 ? $signed(8'sh37) : $signed(_GEN_429); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_431 = 7'h1c == data1Frac_3 ? $signed(8'sh37) : $signed(_GEN_430); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_432 = 7'h1d == data1Frac_3 ? $signed(8'sh37) : $signed(_GEN_431); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_433 = 7'h1e == data1Frac_3 ? $signed(8'sh36) : $signed(_GEN_432); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_434 = 7'h1f == data1Frac_3 ? $signed(8'sh36) : $signed(_GEN_433); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_435 = 7'h20 == data1Frac_3 ? $signed(8'sh36) : $signed(_GEN_434); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_436 = 7'h21 == data1Frac_3 ? $signed(8'sh36) : $signed(_GEN_435); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_437 = 7'h22 == data1Frac_3 ? $signed(8'sh35) : $signed(_GEN_436); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_438 = 7'h23 == data1Frac_3 ? $signed(8'sh35) : $signed(_GEN_437); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_439 = 7'h24 == data1Frac_3 ? $signed(8'sh35) : $signed(_GEN_438); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_440 = 7'h25 == data1Frac_3 ? $signed(8'sh34) : $signed(_GEN_439); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_441 = 7'h26 == data1Frac_3 ? $signed(8'sh34) : $signed(_GEN_440); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_442 = 7'h27 == data1Frac_3 ? $signed(8'sh34) : $signed(_GEN_441); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_443 = 7'h28 == data1Frac_3 ? $signed(8'sh34) : $signed(_GEN_442); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_444 = 7'h29 == data1Frac_3 ? $signed(8'sh33) : $signed(_GEN_443); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_445 = 7'h2a == data1Frac_3 ? $signed(8'sh33) : $signed(_GEN_444); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_446 = 7'h2b == data1Frac_3 ? $signed(8'sh33) : $signed(_GEN_445); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_447 = 7'h2c == data1Frac_3 ? $signed(8'sh32) : $signed(_GEN_446); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_448 = 7'h2d == data1Frac_3 ? $signed(8'sh32) : $signed(_GEN_447); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_449 = 7'h2e == data1Frac_3 ? $signed(8'sh32) : $signed(_GEN_448); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_450 = 7'h2f == data1Frac_3 ? $signed(8'sh32) : $signed(_GEN_449); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_451 = 7'h30 == data1Frac_3 ? $signed(8'sh31) : $signed(_GEN_450); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_452 = 7'h31 == data1Frac_3 ? $signed(8'sh31) : $signed(_GEN_451); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_453 = 7'h32 == data1Frac_3 ? $signed(8'sh31) : $signed(_GEN_452); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_454 = 7'h33 == data1Frac_3 ? $signed(8'sh31) : $signed(_GEN_453); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_455 = 7'h34 == data1Frac_3 ? $signed(8'sh30) : $signed(_GEN_454); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_456 = 7'h35 == data1Frac_3 ? $signed(8'sh30) : $signed(_GEN_455); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_457 = 7'h36 == data1Frac_3 ? $signed(8'sh30) : $signed(_GEN_456); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_458 = 7'h37 == data1Frac_3 ? $signed(8'sh30) : $signed(_GEN_457); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_459 = 7'h38 == data1Frac_3 ? $signed(8'sh2f) : $signed(_GEN_458); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_460 = 7'h39 == data1Frac_3 ? $signed(8'sh2f) : $signed(_GEN_459); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_461 = 7'h3a == data1Frac_3 ? $signed(8'sh2f) : $signed(_GEN_460); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_462 = 7'h3b == data1Frac_3 ? $signed(8'sh2e) : $signed(_GEN_461); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_463 = 7'h3c == data1Frac_3 ? $signed(8'sh2e) : $signed(_GEN_462); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_464 = 7'h3d == data1Frac_3 ? $signed(8'sh2e) : $signed(_GEN_463); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_465 = 7'h3e == data1Frac_3 ? $signed(8'sh2e) : $signed(_GEN_464); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_466 = 7'h3f == data1Frac_3 ? $signed(8'sh2e) : $signed(_GEN_465); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_467 = 7'h40 == data1Frac_3 ? $signed(8'sh2d) : $signed(_GEN_466); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_468 = 7'h41 == data1Frac_3 ? $signed(8'sh2d) : $signed(_GEN_467); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_469 = 7'h42 == data1Frac_3 ? $signed(8'sh2d) : $signed(_GEN_468); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_470 = 7'h43 == data1Frac_3 ? $signed(8'sh2d) : $signed(_GEN_469); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_471 = 7'h44 == data1Frac_3 ? $signed(8'sh2c) : $signed(_GEN_470); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_472 = 7'h45 == data1Frac_3 ? $signed(8'sh2c) : $signed(_GEN_471); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_473 = 7'h46 == data1Frac_3 ? $signed(8'sh2c) : $signed(_GEN_472); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_474 = 7'h47 == data1Frac_3 ? $signed(8'sh2c) : $signed(_GEN_473); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_475 = 7'h48 == data1Frac_3 ? $signed(8'sh2b) : $signed(_GEN_474); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_476 = 7'h49 == data1Frac_3 ? $signed(8'sh2b) : $signed(_GEN_475); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_477 = 7'h4a == data1Frac_3 ? $signed(8'sh2b) : $signed(_GEN_476); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_478 = 7'h4b == data1Frac_3 ? $signed(8'sh2b) : $signed(_GEN_477); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_479 = 7'h4c == data1Frac_3 ? $signed(8'sh2a) : $signed(_GEN_478); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_480 = 7'h4d == data1Frac_3 ? $signed(8'sh2a) : $signed(_GEN_479); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_481 = 7'h4e == data1Frac_3 ? $signed(8'sh2a) : $signed(_GEN_480); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_482 = 7'h4f == data1Frac_3 ? $signed(8'sh2a) : $signed(_GEN_481); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_483 = 7'h50 == data1Frac_3 ? $signed(8'sh29) : $signed(_GEN_482); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_484 = 7'h51 == data1Frac_3 ? $signed(8'sh29) : $signed(_GEN_483); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_485 = 7'h52 == data1Frac_3 ? $signed(8'sh29) : $signed(_GEN_484); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_486 = 7'h53 == data1Frac_3 ? $signed(8'sh29) : $signed(_GEN_485); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_487 = 7'h54 == data1Frac_3 ? $signed(8'sh29) : $signed(_GEN_486); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_488 = 7'h55 == data1Frac_3 ? $signed(8'sh28) : $signed(_GEN_487); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_489 = 7'h56 == data1Frac_3 ? $signed(8'sh28) : $signed(_GEN_488); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_490 = 7'h57 == data1Frac_3 ? $signed(8'sh28) : $signed(_GEN_489); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_491 = 7'h58 == data1Frac_3 ? $signed(8'sh28) : $signed(_GEN_490); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_492 = 7'h59 == data1Frac_3 ? $signed(8'sh28) : $signed(_GEN_491); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_493 = 7'h5a == data1Frac_3 ? $signed(8'sh27) : $signed(_GEN_492); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_494 = 7'h5b == data1Frac_3 ? $signed(8'sh27) : $signed(_GEN_493); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_495 = 7'h5c == data1Frac_3 ? $signed(8'sh27) : $signed(_GEN_494); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_496 = 7'h5d == data1Frac_3 ? $signed(8'sh27) : $signed(_GEN_495); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_497 = 7'h5e == data1Frac_3 ? $signed(8'sh26) : $signed(_GEN_496); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_498 = 7'h5f == data1Frac_3 ? $signed(8'sh26) : $signed(_GEN_497); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_499 = 7'h60 == data1Frac_3 ? $signed(8'sh26) : $signed(_GEN_498); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_500 = 7'h61 == data1Frac_3 ? $signed(8'sh26) : $signed(_GEN_499); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_501 = 7'h62 == data1Frac_3 ? $signed(8'sh26) : $signed(_GEN_500); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_502 = 7'h63 == data1Frac_3 ? $signed(8'sh25) : $signed(_GEN_501); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_503 = 7'h64 == data1Frac_3 ? $signed(8'sh25) : $signed(_GEN_502); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_504 = 7'h65 == data1Frac_3 ? $signed(8'sh25) : $signed(_GEN_503); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_505 = 7'h66 == data1Frac_3 ? $signed(8'sh25) : $signed(_GEN_504); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_506 = 7'h67 == data1Frac_3 ? $signed(8'sh25) : $signed(_GEN_505); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_507 = 7'h68 == data1Frac_3 ? $signed(8'sh24) : $signed(_GEN_506); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_508 = 7'h69 == data1Frac_3 ? $signed(8'sh24) : $signed(_GEN_507); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_509 = 7'h6a == data1Frac_3 ? $signed(8'sh24) : $signed(_GEN_508); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_510 = 7'h6b == data1Frac_3 ? $signed(8'sh24) : $signed(_GEN_509); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_511 = 7'h6c == data1Frac_3 ? $signed(8'sh24) : $signed(_GEN_510); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_512 = 7'h6d == data1Frac_3 ? $signed(8'sh23) : $signed(_GEN_511); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_513 = 7'h6e == data1Frac_3 ? $signed(8'sh23) : $signed(_GEN_512); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_514 = 7'h6f == data1Frac_3 ? $signed(8'sh23) : $signed(_GEN_513); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_515 = 7'h70 == data1Frac_3 ? $signed(8'sh23) : $signed(_GEN_514); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_516 = 7'h71 == data1Frac_3 ? $signed(8'sh23) : $signed(_GEN_515); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_517 = 7'h72 == data1Frac_3 ? $signed(8'sh23) : $signed(_GEN_516); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_518 = 7'h73 == data1Frac_3 ? $signed(8'sh22) : $signed(_GEN_517); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_519 = 7'h74 == data1Frac_3 ? $signed(8'sh22) : $signed(_GEN_518); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_520 = 7'h75 == data1Frac_3 ? $signed(8'sh22) : $signed(_GEN_519); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_521 = 7'h76 == data1Frac_3 ? $signed(8'sh22) : $signed(_GEN_520); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_522 = 7'h77 == data1Frac_3 ? $signed(8'sh22) : $signed(_GEN_521); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_523 = 7'h78 == data1Frac_3 ? $signed(8'sh21) : $signed(_GEN_522); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_524 = 7'h79 == data1Frac_3 ? $signed(8'sh21) : $signed(_GEN_523); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_525 = 7'h7a == data1Frac_3 ? $signed(8'sh21) : $signed(_GEN_524); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_526 = 7'h7b == data1Frac_3 ? $signed(8'sh21) : $signed(_GEN_525); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_527 = 7'h7c == data1Frac_3 ? $signed(8'sh21) : $signed(_GEN_526); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_528 = 7'h7d == data1Frac_3 ? $signed(8'sh21) : $signed(_GEN_527); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_529 = 7'h7e == data1Frac_3 ? $signed(8'sh20) : $signed(_GEN_528); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_530 = 7'h7f == data1Frac_3 ? $signed(8'sh20) : $signed(_GEN_529); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_11 = $signed(_GEN_530) >>> data1Int_3; // @[exponent.scala 38:85]
  reg [7:0] data2_3; // @[Reg.scala 16:16]
  wire [7:0] _GEN_534 = 7'h2 == data1Frac_4 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_535 = 7'h3 == data1Frac_4 ? $signed(8'sh3f) : $signed(_GEN_534); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_536 = 7'h4 == data1Frac_4 ? $signed(8'sh3f) : $signed(_GEN_535); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_537 = 7'h5 == data1Frac_4 ? $signed(8'sh3e) : $signed(_GEN_536); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_538 = 7'h6 == data1Frac_4 ? $signed(8'sh3e) : $signed(_GEN_537); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_539 = 7'h7 == data1Frac_4 ? $signed(8'sh3e) : $signed(_GEN_538); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_540 = 7'h8 == data1Frac_4 ? $signed(8'sh3d) : $signed(_GEN_539); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_541 = 7'h9 == data1Frac_4 ? $signed(8'sh3d) : $signed(_GEN_540); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_542 = 7'ha == data1Frac_4 ? $signed(8'sh3d) : $signed(_GEN_541); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_543 = 7'hb == data1Frac_4 ? $signed(8'sh3c) : $signed(_GEN_542); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_544 = 7'hc == data1Frac_4 ? $signed(8'sh3c) : $signed(_GEN_543); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_545 = 7'hd == data1Frac_4 ? $signed(8'sh3c) : $signed(_GEN_544); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_546 = 7'he == data1Frac_4 ? $signed(8'sh3b) : $signed(_GEN_545); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_547 = 7'hf == data1Frac_4 ? $signed(8'sh3b) : $signed(_GEN_546); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_548 = 7'h10 == data1Frac_4 ? $signed(8'sh3b) : $signed(_GEN_547); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_549 = 7'h11 == data1Frac_4 ? $signed(8'sh3a) : $signed(_GEN_548); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_550 = 7'h12 == data1Frac_4 ? $signed(8'sh3a) : $signed(_GEN_549); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_551 = 7'h13 == data1Frac_4 ? $signed(8'sh3a) : $signed(_GEN_550); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_552 = 7'h14 == data1Frac_4 ? $signed(8'sh39) : $signed(_GEN_551); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_553 = 7'h15 == data1Frac_4 ? $signed(8'sh39) : $signed(_GEN_552); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_554 = 7'h16 == data1Frac_4 ? $signed(8'sh39) : $signed(_GEN_553); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_555 = 7'h17 == data1Frac_4 ? $signed(8'sh39) : $signed(_GEN_554); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_556 = 7'h18 == data1Frac_4 ? $signed(8'sh38) : $signed(_GEN_555); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_557 = 7'h19 == data1Frac_4 ? $signed(8'sh38) : $signed(_GEN_556); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_558 = 7'h1a == data1Frac_4 ? $signed(8'sh38) : $signed(_GEN_557); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_559 = 7'h1b == data1Frac_4 ? $signed(8'sh37) : $signed(_GEN_558); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_560 = 7'h1c == data1Frac_4 ? $signed(8'sh37) : $signed(_GEN_559); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_561 = 7'h1d == data1Frac_4 ? $signed(8'sh37) : $signed(_GEN_560); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_562 = 7'h1e == data1Frac_4 ? $signed(8'sh36) : $signed(_GEN_561); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_563 = 7'h1f == data1Frac_4 ? $signed(8'sh36) : $signed(_GEN_562); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_564 = 7'h20 == data1Frac_4 ? $signed(8'sh36) : $signed(_GEN_563); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_565 = 7'h21 == data1Frac_4 ? $signed(8'sh36) : $signed(_GEN_564); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_566 = 7'h22 == data1Frac_4 ? $signed(8'sh35) : $signed(_GEN_565); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_567 = 7'h23 == data1Frac_4 ? $signed(8'sh35) : $signed(_GEN_566); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_568 = 7'h24 == data1Frac_4 ? $signed(8'sh35) : $signed(_GEN_567); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_569 = 7'h25 == data1Frac_4 ? $signed(8'sh34) : $signed(_GEN_568); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_570 = 7'h26 == data1Frac_4 ? $signed(8'sh34) : $signed(_GEN_569); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_571 = 7'h27 == data1Frac_4 ? $signed(8'sh34) : $signed(_GEN_570); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_572 = 7'h28 == data1Frac_4 ? $signed(8'sh34) : $signed(_GEN_571); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_573 = 7'h29 == data1Frac_4 ? $signed(8'sh33) : $signed(_GEN_572); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_574 = 7'h2a == data1Frac_4 ? $signed(8'sh33) : $signed(_GEN_573); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_575 = 7'h2b == data1Frac_4 ? $signed(8'sh33) : $signed(_GEN_574); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_576 = 7'h2c == data1Frac_4 ? $signed(8'sh32) : $signed(_GEN_575); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_577 = 7'h2d == data1Frac_4 ? $signed(8'sh32) : $signed(_GEN_576); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_578 = 7'h2e == data1Frac_4 ? $signed(8'sh32) : $signed(_GEN_577); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_579 = 7'h2f == data1Frac_4 ? $signed(8'sh32) : $signed(_GEN_578); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_580 = 7'h30 == data1Frac_4 ? $signed(8'sh31) : $signed(_GEN_579); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_581 = 7'h31 == data1Frac_4 ? $signed(8'sh31) : $signed(_GEN_580); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_582 = 7'h32 == data1Frac_4 ? $signed(8'sh31) : $signed(_GEN_581); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_583 = 7'h33 == data1Frac_4 ? $signed(8'sh31) : $signed(_GEN_582); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_584 = 7'h34 == data1Frac_4 ? $signed(8'sh30) : $signed(_GEN_583); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_585 = 7'h35 == data1Frac_4 ? $signed(8'sh30) : $signed(_GEN_584); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_586 = 7'h36 == data1Frac_4 ? $signed(8'sh30) : $signed(_GEN_585); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_587 = 7'h37 == data1Frac_4 ? $signed(8'sh30) : $signed(_GEN_586); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_588 = 7'h38 == data1Frac_4 ? $signed(8'sh2f) : $signed(_GEN_587); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_589 = 7'h39 == data1Frac_4 ? $signed(8'sh2f) : $signed(_GEN_588); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_590 = 7'h3a == data1Frac_4 ? $signed(8'sh2f) : $signed(_GEN_589); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_591 = 7'h3b == data1Frac_4 ? $signed(8'sh2e) : $signed(_GEN_590); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_592 = 7'h3c == data1Frac_4 ? $signed(8'sh2e) : $signed(_GEN_591); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_593 = 7'h3d == data1Frac_4 ? $signed(8'sh2e) : $signed(_GEN_592); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_594 = 7'h3e == data1Frac_4 ? $signed(8'sh2e) : $signed(_GEN_593); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_595 = 7'h3f == data1Frac_4 ? $signed(8'sh2e) : $signed(_GEN_594); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_596 = 7'h40 == data1Frac_4 ? $signed(8'sh2d) : $signed(_GEN_595); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_597 = 7'h41 == data1Frac_4 ? $signed(8'sh2d) : $signed(_GEN_596); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_598 = 7'h42 == data1Frac_4 ? $signed(8'sh2d) : $signed(_GEN_597); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_599 = 7'h43 == data1Frac_4 ? $signed(8'sh2d) : $signed(_GEN_598); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_600 = 7'h44 == data1Frac_4 ? $signed(8'sh2c) : $signed(_GEN_599); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_601 = 7'h45 == data1Frac_4 ? $signed(8'sh2c) : $signed(_GEN_600); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_602 = 7'h46 == data1Frac_4 ? $signed(8'sh2c) : $signed(_GEN_601); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_603 = 7'h47 == data1Frac_4 ? $signed(8'sh2c) : $signed(_GEN_602); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_604 = 7'h48 == data1Frac_4 ? $signed(8'sh2b) : $signed(_GEN_603); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_605 = 7'h49 == data1Frac_4 ? $signed(8'sh2b) : $signed(_GEN_604); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_606 = 7'h4a == data1Frac_4 ? $signed(8'sh2b) : $signed(_GEN_605); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_607 = 7'h4b == data1Frac_4 ? $signed(8'sh2b) : $signed(_GEN_606); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_608 = 7'h4c == data1Frac_4 ? $signed(8'sh2a) : $signed(_GEN_607); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_609 = 7'h4d == data1Frac_4 ? $signed(8'sh2a) : $signed(_GEN_608); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_610 = 7'h4e == data1Frac_4 ? $signed(8'sh2a) : $signed(_GEN_609); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_611 = 7'h4f == data1Frac_4 ? $signed(8'sh2a) : $signed(_GEN_610); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_612 = 7'h50 == data1Frac_4 ? $signed(8'sh29) : $signed(_GEN_611); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_613 = 7'h51 == data1Frac_4 ? $signed(8'sh29) : $signed(_GEN_612); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_614 = 7'h52 == data1Frac_4 ? $signed(8'sh29) : $signed(_GEN_613); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_615 = 7'h53 == data1Frac_4 ? $signed(8'sh29) : $signed(_GEN_614); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_616 = 7'h54 == data1Frac_4 ? $signed(8'sh29) : $signed(_GEN_615); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_617 = 7'h55 == data1Frac_4 ? $signed(8'sh28) : $signed(_GEN_616); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_618 = 7'h56 == data1Frac_4 ? $signed(8'sh28) : $signed(_GEN_617); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_619 = 7'h57 == data1Frac_4 ? $signed(8'sh28) : $signed(_GEN_618); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_620 = 7'h58 == data1Frac_4 ? $signed(8'sh28) : $signed(_GEN_619); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_621 = 7'h59 == data1Frac_4 ? $signed(8'sh28) : $signed(_GEN_620); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_622 = 7'h5a == data1Frac_4 ? $signed(8'sh27) : $signed(_GEN_621); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_623 = 7'h5b == data1Frac_4 ? $signed(8'sh27) : $signed(_GEN_622); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_624 = 7'h5c == data1Frac_4 ? $signed(8'sh27) : $signed(_GEN_623); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_625 = 7'h5d == data1Frac_4 ? $signed(8'sh27) : $signed(_GEN_624); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_626 = 7'h5e == data1Frac_4 ? $signed(8'sh26) : $signed(_GEN_625); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_627 = 7'h5f == data1Frac_4 ? $signed(8'sh26) : $signed(_GEN_626); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_628 = 7'h60 == data1Frac_4 ? $signed(8'sh26) : $signed(_GEN_627); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_629 = 7'h61 == data1Frac_4 ? $signed(8'sh26) : $signed(_GEN_628); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_630 = 7'h62 == data1Frac_4 ? $signed(8'sh26) : $signed(_GEN_629); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_631 = 7'h63 == data1Frac_4 ? $signed(8'sh25) : $signed(_GEN_630); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_632 = 7'h64 == data1Frac_4 ? $signed(8'sh25) : $signed(_GEN_631); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_633 = 7'h65 == data1Frac_4 ? $signed(8'sh25) : $signed(_GEN_632); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_634 = 7'h66 == data1Frac_4 ? $signed(8'sh25) : $signed(_GEN_633); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_635 = 7'h67 == data1Frac_4 ? $signed(8'sh25) : $signed(_GEN_634); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_636 = 7'h68 == data1Frac_4 ? $signed(8'sh24) : $signed(_GEN_635); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_637 = 7'h69 == data1Frac_4 ? $signed(8'sh24) : $signed(_GEN_636); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_638 = 7'h6a == data1Frac_4 ? $signed(8'sh24) : $signed(_GEN_637); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_639 = 7'h6b == data1Frac_4 ? $signed(8'sh24) : $signed(_GEN_638); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_640 = 7'h6c == data1Frac_4 ? $signed(8'sh24) : $signed(_GEN_639); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_641 = 7'h6d == data1Frac_4 ? $signed(8'sh23) : $signed(_GEN_640); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_642 = 7'h6e == data1Frac_4 ? $signed(8'sh23) : $signed(_GEN_641); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_643 = 7'h6f == data1Frac_4 ? $signed(8'sh23) : $signed(_GEN_642); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_644 = 7'h70 == data1Frac_4 ? $signed(8'sh23) : $signed(_GEN_643); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_645 = 7'h71 == data1Frac_4 ? $signed(8'sh23) : $signed(_GEN_644); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_646 = 7'h72 == data1Frac_4 ? $signed(8'sh23) : $signed(_GEN_645); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_647 = 7'h73 == data1Frac_4 ? $signed(8'sh22) : $signed(_GEN_646); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_648 = 7'h74 == data1Frac_4 ? $signed(8'sh22) : $signed(_GEN_647); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_649 = 7'h75 == data1Frac_4 ? $signed(8'sh22) : $signed(_GEN_648); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_650 = 7'h76 == data1Frac_4 ? $signed(8'sh22) : $signed(_GEN_649); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_651 = 7'h77 == data1Frac_4 ? $signed(8'sh22) : $signed(_GEN_650); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_652 = 7'h78 == data1Frac_4 ? $signed(8'sh21) : $signed(_GEN_651); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_653 = 7'h79 == data1Frac_4 ? $signed(8'sh21) : $signed(_GEN_652); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_654 = 7'h7a == data1Frac_4 ? $signed(8'sh21) : $signed(_GEN_653); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_655 = 7'h7b == data1Frac_4 ? $signed(8'sh21) : $signed(_GEN_654); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_656 = 7'h7c == data1Frac_4 ? $signed(8'sh21) : $signed(_GEN_655); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_657 = 7'h7d == data1Frac_4 ? $signed(8'sh21) : $signed(_GEN_656); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_658 = 7'h7e == data1Frac_4 ? $signed(8'sh20) : $signed(_GEN_657); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_659 = 7'h7f == data1Frac_4 ? $signed(8'sh20) : $signed(_GEN_658); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_14 = $signed(_GEN_659) >>> data1Int_4; // @[exponent.scala 38:85]
  reg [7:0] data2_4; // @[Reg.scala 16:16]
  wire [7:0] _GEN_663 = 7'h2 == data1Frac_5 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_664 = 7'h3 == data1Frac_5 ? $signed(8'sh3f) : $signed(_GEN_663); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_665 = 7'h4 == data1Frac_5 ? $signed(8'sh3f) : $signed(_GEN_664); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_666 = 7'h5 == data1Frac_5 ? $signed(8'sh3e) : $signed(_GEN_665); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_667 = 7'h6 == data1Frac_5 ? $signed(8'sh3e) : $signed(_GEN_666); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_668 = 7'h7 == data1Frac_5 ? $signed(8'sh3e) : $signed(_GEN_667); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_669 = 7'h8 == data1Frac_5 ? $signed(8'sh3d) : $signed(_GEN_668); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_670 = 7'h9 == data1Frac_5 ? $signed(8'sh3d) : $signed(_GEN_669); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_671 = 7'ha == data1Frac_5 ? $signed(8'sh3d) : $signed(_GEN_670); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_672 = 7'hb == data1Frac_5 ? $signed(8'sh3c) : $signed(_GEN_671); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_673 = 7'hc == data1Frac_5 ? $signed(8'sh3c) : $signed(_GEN_672); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_674 = 7'hd == data1Frac_5 ? $signed(8'sh3c) : $signed(_GEN_673); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_675 = 7'he == data1Frac_5 ? $signed(8'sh3b) : $signed(_GEN_674); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_676 = 7'hf == data1Frac_5 ? $signed(8'sh3b) : $signed(_GEN_675); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_677 = 7'h10 == data1Frac_5 ? $signed(8'sh3b) : $signed(_GEN_676); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_678 = 7'h11 == data1Frac_5 ? $signed(8'sh3a) : $signed(_GEN_677); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_679 = 7'h12 == data1Frac_5 ? $signed(8'sh3a) : $signed(_GEN_678); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_680 = 7'h13 == data1Frac_5 ? $signed(8'sh3a) : $signed(_GEN_679); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_681 = 7'h14 == data1Frac_5 ? $signed(8'sh39) : $signed(_GEN_680); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_682 = 7'h15 == data1Frac_5 ? $signed(8'sh39) : $signed(_GEN_681); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_683 = 7'h16 == data1Frac_5 ? $signed(8'sh39) : $signed(_GEN_682); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_684 = 7'h17 == data1Frac_5 ? $signed(8'sh39) : $signed(_GEN_683); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_685 = 7'h18 == data1Frac_5 ? $signed(8'sh38) : $signed(_GEN_684); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_686 = 7'h19 == data1Frac_5 ? $signed(8'sh38) : $signed(_GEN_685); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_687 = 7'h1a == data1Frac_5 ? $signed(8'sh38) : $signed(_GEN_686); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_688 = 7'h1b == data1Frac_5 ? $signed(8'sh37) : $signed(_GEN_687); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_689 = 7'h1c == data1Frac_5 ? $signed(8'sh37) : $signed(_GEN_688); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_690 = 7'h1d == data1Frac_5 ? $signed(8'sh37) : $signed(_GEN_689); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_691 = 7'h1e == data1Frac_5 ? $signed(8'sh36) : $signed(_GEN_690); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_692 = 7'h1f == data1Frac_5 ? $signed(8'sh36) : $signed(_GEN_691); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_693 = 7'h20 == data1Frac_5 ? $signed(8'sh36) : $signed(_GEN_692); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_694 = 7'h21 == data1Frac_5 ? $signed(8'sh36) : $signed(_GEN_693); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_695 = 7'h22 == data1Frac_5 ? $signed(8'sh35) : $signed(_GEN_694); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_696 = 7'h23 == data1Frac_5 ? $signed(8'sh35) : $signed(_GEN_695); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_697 = 7'h24 == data1Frac_5 ? $signed(8'sh35) : $signed(_GEN_696); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_698 = 7'h25 == data1Frac_5 ? $signed(8'sh34) : $signed(_GEN_697); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_699 = 7'h26 == data1Frac_5 ? $signed(8'sh34) : $signed(_GEN_698); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_700 = 7'h27 == data1Frac_5 ? $signed(8'sh34) : $signed(_GEN_699); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_701 = 7'h28 == data1Frac_5 ? $signed(8'sh34) : $signed(_GEN_700); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_702 = 7'h29 == data1Frac_5 ? $signed(8'sh33) : $signed(_GEN_701); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_703 = 7'h2a == data1Frac_5 ? $signed(8'sh33) : $signed(_GEN_702); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_704 = 7'h2b == data1Frac_5 ? $signed(8'sh33) : $signed(_GEN_703); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_705 = 7'h2c == data1Frac_5 ? $signed(8'sh32) : $signed(_GEN_704); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_706 = 7'h2d == data1Frac_5 ? $signed(8'sh32) : $signed(_GEN_705); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_707 = 7'h2e == data1Frac_5 ? $signed(8'sh32) : $signed(_GEN_706); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_708 = 7'h2f == data1Frac_5 ? $signed(8'sh32) : $signed(_GEN_707); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_709 = 7'h30 == data1Frac_5 ? $signed(8'sh31) : $signed(_GEN_708); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_710 = 7'h31 == data1Frac_5 ? $signed(8'sh31) : $signed(_GEN_709); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_711 = 7'h32 == data1Frac_5 ? $signed(8'sh31) : $signed(_GEN_710); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_712 = 7'h33 == data1Frac_5 ? $signed(8'sh31) : $signed(_GEN_711); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_713 = 7'h34 == data1Frac_5 ? $signed(8'sh30) : $signed(_GEN_712); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_714 = 7'h35 == data1Frac_5 ? $signed(8'sh30) : $signed(_GEN_713); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_715 = 7'h36 == data1Frac_5 ? $signed(8'sh30) : $signed(_GEN_714); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_716 = 7'h37 == data1Frac_5 ? $signed(8'sh30) : $signed(_GEN_715); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_717 = 7'h38 == data1Frac_5 ? $signed(8'sh2f) : $signed(_GEN_716); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_718 = 7'h39 == data1Frac_5 ? $signed(8'sh2f) : $signed(_GEN_717); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_719 = 7'h3a == data1Frac_5 ? $signed(8'sh2f) : $signed(_GEN_718); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_720 = 7'h3b == data1Frac_5 ? $signed(8'sh2e) : $signed(_GEN_719); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_721 = 7'h3c == data1Frac_5 ? $signed(8'sh2e) : $signed(_GEN_720); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_722 = 7'h3d == data1Frac_5 ? $signed(8'sh2e) : $signed(_GEN_721); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_723 = 7'h3e == data1Frac_5 ? $signed(8'sh2e) : $signed(_GEN_722); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_724 = 7'h3f == data1Frac_5 ? $signed(8'sh2e) : $signed(_GEN_723); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_725 = 7'h40 == data1Frac_5 ? $signed(8'sh2d) : $signed(_GEN_724); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_726 = 7'h41 == data1Frac_5 ? $signed(8'sh2d) : $signed(_GEN_725); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_727 = 7'h42 == data1Frac_5 ? $signed(8'sh2d) : $signed(_GEN_726); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_728 = 7'h43 == data1Frac_5 ? $signed(8'sh2d) : $signed(_GEN_727); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_729 = 7'h44 == data1Frac_5 ? $signed(8'sh2c) : $signed(_GEN_728); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_730 = 7'h45 == data1Frac_5 ? $signed(8'sh2c) : $signed(_GEN_729); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_731 = 7'h46 == data1Frac_5 ? $signed(8'sh2c) : $signed(_GEN_730); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_732 = 7'h47 == data1Frac_5 ? $signed(8'sh2c) : $signed(_GEN_731); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_733 = 7'h48 == data1Frac_5 ? $signed(8'sh2b) : $signed(_GEN_732); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_734 = 7'h49 == data1Frac_5 ? $signed(8'sh2b) : $signed(_GEN_733); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_735 = 7'h4a == data1Frac_5 ? $signed(8'sh2b) : $signed(_GEN_734); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_736 = 7'h4b == data1Frac_5 ? $signed(8'sh2b) : $signed(_GEN_735); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_737 = 7'h4c == data1Frac_5 ? $signed(8'sh2a) : $signed(_GEN_736); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_738 = 7'h4d == data1Frac_5 ? $signed(8'sh2a) : $signed(_GEN_737); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_739 = 7'h4e == data1Frac_5 ? $signed(8'sh2a) : $signed(_GEN_738); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_740 = 7'h4f == data1Frac_5 ? $signed(8'sh2a) : $signed(_GEN_739); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_741 = 7'h50 == data1Frac_5 ? $signed(8'sh29) : $signed(_GEN_740); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_742 = 7'h51 == data1Frac_5 ? $signed(8'sh29) : $signed(_GEN_741); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_743 = 7'h52 == data1Frac_5 ? $signed(8'sh29) : $signed(_GEN_742); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_744 = 7'h53 == data1Frac_5 ? $signed(8'sh29) : $signed(_GEN_743); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_745 = 7'h54 == data1Frac_5 ? $signed(8'sh29) : $signed(_GEN_744); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_746 = 7'h55 == data1Frac_5 ? $signed(8'sh28) : $signed(_GEN_745); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_747 = 7'h56 == data1Frac_5 ? $signed(8'sh28) : $signed(_GEN_746); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_748 = 7'h57 == data1Frac_5 ? $signed(8'sh28) : $signed(_GEN_747); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_749 = 7'h58 == data1Frac_5 ? $signed(8'sh28) : $signed(_GEN_748); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_750 = 7'h59 == data1Frac_5 ? $signed(8'sh28) : $signed(_GEN_749); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_751 = 7'h5a == data1Frac_5 ? $signed(8'sh27) : $signed(_GEN_750); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_752 = 7'h5b == data1Frac_5 ? $signed(8'sh27) : $signed(_GEN_751); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_753 = 7'h5c == data1Frac_5 ? $signed(8'sh27) : $signed(_GEN_752); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_754 = 7'h5d == data1Frac_5 ? $signed(8'sh27) : $signed(_GEN_753); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_755 = 7'h5e == data1Frac_5 ? $signed(8'sh26) : $signed(_GEN_754); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_756 = 7'h5f == data1Frac_5 ? $signed(8'sh26) : $signed(_GEN_755); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_757 = 7'h60 == data1Frac_5 ? $signed(8'sh26) : $signed(_GEN_756); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_758 = 7'h61 == data1Frac_5 ? $signed(8'sh26) : $signed(_GEN_757); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_759 = 7'h62 == data1Frac_5 ? $signed(8'sh26) : $signed(_GEN_758); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_760 = 7'h63 == data1Frac_5 ? $signed(8'sh25) : $signed(_GEN_759); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_761 = 7'h64 == data1Frac_5 ? $signed(8'sh25) : $signed(_GEN_760); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_762 = 7'h65 == data1Frac_5 ? $signed(8'sh25) : $signed(_GEN_761); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_763 = 7'h66 == data1Frac_5 ? $signed(8'sh25) : $signed(_GEN_762); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_764 = 7'h67 == data1Frac_5 ? $signed(8'sh25) : $signed(_GEN_763); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_765 = 7'h68 == data1Frac_5 ? $signed(8'sh24) : $signed(_GEN_764); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_766 = 7'h69 == data1Frac_5 ? $signed(8'sh24) : $signed(_GEN_765); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_767 = 7'h6a == data1Frac_5 ? $signed(8'sh24) : $signed(_GEN_766); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_768 = 7'h6b == data1Frac_5 ? $signed(8'sh24) : $signed(_GEN_767); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_769 = 7'h6c == data1Frac_5 ? $signed(8'sh24) : $signed(_GEN_768); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_770 = 7'h6d == data1Frac_5 ? $signed(8'sh23) : $signed(_GEN_769); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_771 = 7'h6e == data1Frac_5 ? $signed(8'sh23) : $signed(_GEN_770); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_772 = 7'h6f == data1Frac_5 ? $signed(8'sh23) : $signed(_GEN_771); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_773 = 7'h70 == data1Frac_5 ? $signed(8'sh23) : $signed(_GEN_772); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_774 = 7'h71 == data1Frac_5 ? $signed(8'sh23) : $signed(_GEN_773); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_775 = 7'h72 == data1Frac_5 ? $signed(8'sh23) : $signed(_GEN_774); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_776 = 7'h73 == data1Frac_5 ? $signed(8'sh22) : $signed(_GEN_775); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_777 = 7'h74 == data1Frac_5 ? $signed(8'sh22) : $signed(_GEN_776); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_778 = 7'h75 == data1Frac_5 ? $signed(8'sh22) : $signed(_GEN_777); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_779 = 7'h76 == data1Frac_5 ? $signed(8'sh22) : $signed(_GEN_778); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_780 = 7'h77 == data1Frac_5 ? $signed(8'sh22) : $signed(_GEN_779); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_781 = 7'h78 == data1Frac_5 ? $signed(8'sh21) : $signed(_GEN_780); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_782 = 7'h79 == data1Frac_5 ? $signed(8'sh21) : $signed(_GEN_781); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_783 = 7'h7a == data1Frac_5 ? $signed(8'sh21) : $signed(_GEN_782); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_784 = 7'h7b == data1Frac_5 ? $signed(8'sh21) : $signed(_GEN_783); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_785 = 7'h7c == data1Frac_5 ? $signed(8'sh21) : $signed(_GEN_784); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_786 = 7'h7d == data1Frac_5 ? $signed(8'sh21) : $signed(_GEN_785); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_787 = 7'h7e == data1Frac_5 ? $signed(8'sh20) : $signed(_GEN_786); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_788 = 7'h7f == data1Frac_5 ? $signed(8'sh20) : $signed(_GEN_787); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_17 = $signed(_GEN_788) >>> data1Int_5; // @[exponent.scala 38:85]
  reg [7:0] data2_5; // @[Reg.scala 16:16]
  wire [7:0] _GEN_792 = 7'h2 == data1Frac_6 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_793 = 7'h3 == data1Frac_6 ? $signed(8'sh3f) : $signed(_GEN_792); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_794 = 7'h4 == data1Frac_6 ? $signed(8'sh3f) : $signed(_GEN_793); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_795 = 7'h5 == data1Frac_6 ? $signed(8'sh3e) : $signed(_GEN_794); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_796 = 7'h6 == data1Frac_6 ? $signed(8'sh3e) : $signed(_GEN_795); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_797 = 7'h7 == data1Frac_6 ? $signed(8'sh3e) : $signed(_GEN_796); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_798 = 7'h8 == data1Frac_6 ? $signed(8'sh3d) : $signed(_GEN_797); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_799 = 7'h9 == data1Frac_6 ? $signed(8'sh3d) : $signed(_GEN_798); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_800 = 7'ha == data1Frac_6 ? $signed(8'sh3d) : $signed(_GEN_799); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_801 = 7'hb == data1Frac_6 ? $signed(8'sh3c) : $signed(_GEN_800); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_802 = 7'hc == data1Frac_6 ? $signed(8'sh3c) : $signed(_GEN_801); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_803 = 7'hd == data1Frac_6 ? $signed(8'sh3c) : $signed(_GEN_802); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_804 = 7'he == data1Frac_6 ? $signed(8'sh3b) : $signed(_GEN_803); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_805 = 7'hf == data1Frac_6 ? $signed(8'sh3b) : $signed(_GEN_804); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_806 = 7'h10 == data1Frac_6 ? $signed(8'sh3b) : $signed(_GEN_805); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_807 = 7'h11 == data1Frac_6 ? $signed(8'sh3a) : $signed(_GEN_806); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_808 = 7'h12 == data1Frac_6 ? $signed(8'sh3a) : $signed(_GEN_807); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_809 = 7'h13 == data1Frac_6 ? $signed(8'sh3a) : $signed(_GEN_808); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_810 = 7'h14 == data1Frac_6 ? $signed(8'sh39) : $signed(_GEN_809); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_811 = 7'h15 == data1Frac_6 ? $signed(8'sh39) : $signed(_GEN_810); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_812 = 7'h16 == data1Frac_6 ? $signed(8'sh39) : $signed(_GEN_811); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_813 = 7'h17 == data1Frac_6 ? $signed(8'sh39) : $signed(_GEN_812); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_814 = 7'h18 == data1Frac_6 ? $signed(8'sh38) : $signed(_GEN_813); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_815 = 7'h19 == data1Frac_6 ? $signed(8'sh38) : $signed(_GEN_814); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_816 = 7'h1a == data1Frac_6 ? $signed(8'sh38) : $signed(_GEN_815); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_817 = 7'h1b == data1Frac_6 ? $signed(8'sh37) : $signed(_GEN_816); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_818 = 7'h1c == data1Frac_6 ? $signed(8'sh37) : $signed(_GEN_817); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_819 = 7'h1d == data1Frac_6 ? $signed(8'sh37) : $signed(_GEN_818); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_820 = 7'h1e == data1Frac_6 ? $signed(8'sh36) : $signed(_GEN_819); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_821 = 7'h1f == data1Frac_6 ? $signed(8'sh36) : $signed(_GEN_820); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_822 = 7'h20 == data1Frac_6 ? $signed(8'sh36) : $signed(_GEN_821); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_823 = 7'h21 == data1Frac_6 ? $signed(8'sh36) : $signed(_GEN_822); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_824 = 7'h22 == data1Frac_6 ? $signed(8'sh35) : $signed(_GEN_823); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_825 = 7'h23 == data1Frac_6 ? $signed(8'sh35) : $signed(_GEN_824); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_826 = 7'h24 == data1Frac_6 ? $signed(8'sh35) : $signed(_GEN_825); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_827 = 7'h25 == data1Frac_6 ? $signed(8'sh34) : $signed(_GEN_826); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_828 = 7'h26 == data1Frac_6 ? $signed(8'sh34) : $signed(_GEN_827); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_829 = 7'h27 == data1Frac_6 ? $signed(8'sh34) : $signed(_GEN_828); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_830 = 7'h28 == data1Frac_6 ? $signed(8'sh34) : $signed(_GEN_829); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_831 = 7'h29 == data1Frac_6 ? $signed(8'sh33) : $signed(_GEN_830); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_832 = 7'h2a == data1Frac_6 ? $signed(8'sh33) : $signed(_GEN_831); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_833 = 7'h2b == data1Frac_6 ? $signed(8'sh33) : $signed(_GEN_832); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_834 = 7'h2c == data1Frac_6 ? $signed(8'sh32) : $signed(_GEN_833); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_835 = 7'h2d == data1Frac_6 ? $signed(8'sh32) : $signed(_GEN_834); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_836 = 7'h2e == data1Frac_6 ? $signed(8'sh32) : $signed(_GEN_835); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_837 = 7'h2f == data1Frac_6 ? $signed(8'sh32) : $signed(_GEN_836); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_838 = 7'h30 == data1Frac_6 ? $signed(8'sh31) : $signed(_GEN_837); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_839 = 7'h31 == data1Frac_6 ? $signed(8'sh31) : $signed(_GEN_838); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_840 = 7'h32 == data1Frac_6 ? $signed(8'sh31) : $signed(_GEN_839); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_841 = 7'h33 == data1Frac_6 ? $signed(8'sh31) : $signed(_GEN_840); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_842 = 7'h34 == data1Frac_6 ? $signed(8'sh30) : $signed(_GEN_841); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_843 = 7'h35 == data1Frac_6 ? $signed(8'sh30) : $signed(_GEN_842); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_844 = 7'h36 == data1Frac_6 ? $signed(8'sh30) : $signed(_GEN_843); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_845 = 7'h37 == data1Frac_6 ? $signed(8'sh30) : $signed(_GEN_844); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_846 = 7'h38 == data1Frac_6 ? $signed(8'sh2f) : $signed(_GEN_845); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_847 = 7'h39 == data1Frac_6 ? $signed(8'sh2f) : $signed(_GEN_846); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_848 = 7'h3a == data1Frac_6 ? $signed(8'sh2f) : $signed(_GEN_847); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_849 = 7'h3b == data1Frac_6 ? $signed(8'sh2e) : $signed(_GEN_848); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_850 = 7'h3c == data1Frac_6 ? $signed(8'sh2e) : $signed(_GEN_849); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_851 = 7'h3d == data1Frac_6 ? $signed(8'sh2e) : $signed(_GEN_850); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_852 = 7'h3e == data1Frac_6 ? $signed(8'sh2e) : $signed(_GEN_851); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_853 = 7'h3f == data1Frac_6 ? $signed(8'sh2e) : $signed(_GEN_852); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_854 = 7'h40 == data1Frac_6 ? $signed(8'sh2d) : $signed(_GEN_853); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_855 = 7'h41 == data1Frac_6 ? $signed(8'sh2d) : $signed(_GEN_854); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_856 = 7'h42 == data1Frac_6 ? $signed(8'sh2d) : $signed(_GEN_855); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_857 = 7'h43 == data1Frac_6 ? $signed(8'sh2d) : $signed(_GEN_856); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_858 = 7'h44 == data1Frac_6 ? $signed(8'sh2c) : $signed(_GEN_857); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_859 = 7'h45 == data1Frac_6 ? $signed(8'sh2c) : $signed(_GEN_858); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_860 = 7'h46 == data1Frac_6 ? $signed(8'sh2c) : $signed(_GEN_859); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_861 = 7'h47 == data1Frac_6 ? $signed(8'sh2c) : $signed(_GEN_860); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_862 = 7'h48 == data1Frac_6 ? $signed(8'sh2b) : $signed(_GEN_861); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_863 = 7'h49 == data1Frac_6 ? $signed(8'sh2b) : $signed(_GEN_862); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_864 = 7'h4a == data1Frac_6 ? $signed(8'sh2b) : $signed(_GEN_863); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_865 = 7'h4b == data1Frac_6 ? $signed(8'sh2b) : $signed(_GEN_864); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_866 = 7'h4c == data1Frac_6 ? $signed(8'sh2a) : $signed(_GEN_865); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_867 = 7'h4d == data1Frac_6 ? $signed(8'sh2a) : $signed(_GEN_866); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_868 = 7'h4e == data1Frac_6 ? $signed(8'sh2a) : $signed(_GEN_867); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_869 = 7'h4f == data1Frac_6 ? $signed(8'sh2a) : $signed(_GEN_868); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_870 = 7'h50 == data1Frac_6 ? $signed(8'sh29) : $signed(_GEN_869); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_871 = 7'h51 == data1Frac_6 ? $signed(8'sh29) : $signed(_GEN_870); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_872 = 7'h52 == data1Frac_6 ? $signed(8'sh29) : $signed(_GEN_871); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_873 = 7'h53 == data1Frac_6 ? $signed(8'sh29) : $signed(_GEN_872); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_874 = 7'h54 == data1Frac_6 ? $signed(8'sh29) : $signed(_GEN_873); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_875 = 7'h55 == data1Frac_6 ? $signed(8'sh28) : $signed(_GEN_874); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_876 = 7'h56 == data1Frac_6 ? $signed(8'sh28) : $signed(_GEN_875); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_877 = 7'h57 == data1Frac_6 ? $signed(8'sh28) : $signed(_GEN_876); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_878 = 7'h58 == data1Frac_6 ? $signed(8'sh28) : $signed(_GEN_877); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_879 = 7'h59 == data1Frac_6 ? $signed(8'sh28) : $signed(_GEN_878); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_880 = 7'h5a == data1Frac_6 ? $signed(8'sh27) : $signed(_GEN_879); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_881 = 7'h5b == data1Frac_6 ? $signed(8'sh27) : $signed(_GEN_880); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_882 = 7'h5c == data1Frac_6 ? $signed(8'sh27) : $signed(_GEN_881); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_883 = 7'h5d == data1Frac_6 ? $signed(8'sh27) : $signed(_GEN_882); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_884 = 7'h5e == data1Frac_6 ? $signed(8'sh26) : $signed(_GEN_883); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_885 = 7'h5f == data1Frac_6 ? $signed(8'sh26) : $signed(_GEN_884); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_886 = 7'h60 == data1Frac_6 ? $signed(8'sh26) : $signed(_GEN_885); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_887 = 7'h61 == data1Frac_6 ? $signed(8'sh26) : $signed(_GEN_886); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_888 = 7'h62 == data1Frac_6 ? $signed(8'sh26) : $signed(_GEN_887); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_889 = 7'h63 == data1Frac_6 ? $signed(8'sh25) : $signed(_GEN_888); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_890 = 7'h64 == data1Frac_6 ? $signed(8'sh25) : $signed(_GEN_889); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_891 = 7'h65 == data1Frac_6 ? $signed(8'sh25) : $signed(_GEN_890); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_892 = 7'h66 == data1Frac_6 ? $signed(8'sh25) : $signed(_GEN_891); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_893 = 7'h67 == data1Frac_6 ? $signed(8'sh25) : $signed(_GEN_892); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_894 = 7'h68 == data1Frac_6 ? $signed(8'sh24) : $signed(_GEN_893); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_895 = 7'h69 == data1Frac_6 ? $signed(8'sh24) : $signed(_GEN_894); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_896 = 7'h6a == data1Frac_6 ? $signed(8'sh24) : $signed(_GEN_895); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_897 = 7'h6b == data1Frac_6 ? $signed(8'sh24) : $signed(_GEN_896); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_898 = 7'h6c == data1Frac_6 ? $signed(8'sh24) : $signed(_GEN_897); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_899 = 7'h6d == data1Frac_6 ? $signed(8'sh23) : $signed(_GEN_898); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_900 = 7'h6e == data1Frac_6 ? $signed(8'sh23) : $signed(_GEN_899); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_901 = 7'h6f == data1Frac_6 ? $signed(8'sh23) : $signed(_GEN_900); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_902 = 7'h70 == data1Frac_6 ? $signed(8'sh23) : $signed(_GEN_901); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_903 = 7'h71 == data1Frac_6 ? $signed(8'sh23) : $signed(_GEN_902); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_904 = 7'h72 == data1Frac_6 ? $signed(8'sh23) : $signed(_GEN_903); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_905 = 7'h73 == data1Frac_6 ? $signed(8'sh22) : $signed(_GEN_904); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_906 = 7'h74 == data1Frac_6 ? $signed(8'sh22) : $signed(_GEN_905); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_907 = 7'h75 == data1Frac_6 ? $signed(8'sh22) : $signed(_GEN_906); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_908 = 7'h76 == data1Frac_6 ? $signed(8'sh22) : $signed(_GEN_907); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_909 = 7'h77 == data1Frac_6 ? $signed(8'sh22) : $signed(_GEN_908); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_910 = 7'h78 == data1Frac_6 ? $signed(8'sh21) : $signed(_GEN_909); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_911 = 7'h79 == data1Frac_6 ? $signed(8'sh21) : $signed(_GEN_910); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_912 = 7'h7a == data1Frac_6 ? $signed(8'sh21) : $signed(_GEN_911); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_913 = 7'h7b == data1Frac_6 ? $signed(8'sh21) : $signed(_GEN_912); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_914 = 7'h7c == data1Frac_6 ? $signed(8'sh21) : $signed(_GEN_913); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_915 = 7'h7d == data1Frac_6 ? $signed(8'sh21) : $signed(_GEN_914); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_916 = 7'h7e == data1Frac_6 ? $signed(8'sh20) : $signed(_GEN_915); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_917 = 7'h7f == data1Frac_6 ? $signed(8'sh20) : $signed(_GEN_916); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_20 = $signed(_GEN_917) >>> data1Int_6; // @[exponent.scala 38:85]
  reg [7:0] data2_6; // @[Reg.scala 16:16]
  wire [7:0] _GEN_921 = 7'h2 == data1Frac_7 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_922 = 7'h3 == data1Frac_7 ? $signed(8'sh3f) : $signed(_GEN_921); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_923 = 7'h4 == data1Frac_7 ? $signed(8'sh3f) : $signed(_GEN_922); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_924 = 7'h5 == data1Frac_7 ? $signed(8'sh3e) : $signed(_GEN_923); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_925 = 7'h6 == data1Frac_7 ? $signed(8'sh3e) : $signed(_GEN_924); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_926 = 7'h7 == data1Frac_7 ? $signed(8'sh3e) : $signed(_GEN_925); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_927 = 7'h8 == data1Frac_7 ? $signed(8'sh3d) : $signed(_GEN_926); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_928 = 7'h9 == data1Frac_7 ? $signed(8'sh3d) : $signed(_GEN_927); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_929 = 7'ha == data1Frac_7 ? $signed(8'sh3d) : $signed(_GEN_928); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_930 = 7'hb == data1Frac_7 ? $signed(8'sh3c) : $signed(_GEN_929); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_931 = 7'hc == data1Frac_7 ? $signed(8'sh3c) : $signed(_GEN_930); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_932 = 7'hd == data1Frac_7 ? $signed(8'sh3c) : $signed(_GEN_931); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_933 = 7'he == data1Frac_7 ? $signed(8'sh3b) : $signed(_GEN_932); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_934 = 7'hf == data1Frac_7 ? $signed(8'sh3b) : $signed(_GEN_933); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_935 = 7'h10 == data1Frac_7 ? $signed(8'sh3b) : $signed(_GEN_934); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_936 = 7'h11 == data1Frac_7 ? $signed(8'sh3a) : $signed(_GEN_935); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_937 = 7'h12 == data1Frac_7 ? $signed(8'sh3a) : $signed(_GEN_936); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_938 = 7'h13 == data1Frac_7 ? $signed(8'sh3a) : $signed(_GEN_937); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_939 = 7'h14 == data1Frac_7 ? $signed(8'sh39) : $signed(_GEN_938); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_940 = 7'h15 == data1Frac_7 ? $signed(8'sh39) : $signed(_GEN_939); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_941 = 7'h16 == data1Frac_7 ? $signed(8'sh39) : $signed(_GEN_940); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_942 = 7'h17 == data1Frac_7 ? $signed(8'sh39) : $signed(_GEN_941); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_943 = 7'h18 == data1Frac_7 ? $signed(8'sh38) : $signed(_GEN_942); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_944 = 7'h19 == data1Frac_7 ? $signed(8'sh38) : $signed(_GEN_943); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_945 = 7'h1a == data1Frac_7 ? $signed(8'sh38) : $signed(_GEN_944); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_946 = 7'h1b == data1Frac_7 ? $signed(8'sh37) : $signed(_GEN_945); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_947 = 7'h1c == data1Frac_7 ? $signed(8'sh37) : $signed(_GEN_946); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_948 = 7'h1d == data1Frac_7 ? $signed(8'sh37) : $signed(_GEN_947); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_949 = 7'h1e == data1Frac_7 ? $signed(8'sh36) : $signed(_GEN_948); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_950 = 7'h1f == data1Frac_7 ? $signed(8'sh36) : $signed(_GEN_949); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_951 = 7'h20 == data1Frac_7 ? $signed(8'sh36) : $signed(_GEN_950); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_952 = 7'h21 == data1Frac_7 ? $signed(8'sh36) : $signed(_GEN_951); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_953 = 7'h22 == data1Frac_7 ? $signed(8'sh35) : $signed(_GEN_952); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_954 = 7'h23 == data1Frac_7 ? $signed(8'sh35) : $signed(_GEN_953); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_955 = 7'h24 == data1Frac_7 ? $signed(8'sh35) : $signed(_GEN_954); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_956 = 7'h25 == data1Frac_7 ? $signed(8'sh34) : $signed(_GEN_955); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_957 = 7'h26 == data1Frac_7 ? $signed(8'sh34) : $signed(_GEN_956); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_958 = 7'h27 == data1Frac_7 ? $signed(8'sh34) : $signed(_GEN_957); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_959 = 7'h28 == data1Frac_7 ? $signed(8'sh34) : $signed(_GEN_958); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_960 = 7'h29 == data1Frac_7 ? $signed(8'sh33) : $signed(_GEN_959); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_961 = 7'h2a == data1Frac_7 ? $signed(8'sh33) : $signed(_GEN_960); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_962 = 7'h2b == data1Frac_7 ? $signed(8'sh33) : $signed(_GEN_961); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_963 = 7'h2c == data1Frac_7 ? $signed(8'sh32) : $signed(_GEN_962); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_964 = 7'h2d == data1Frac_7 ? $signed(8'sh32) : $signed(_GEN_963); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_965 = 7'h2e == data1Frac_7 ? $signed(8'sh32) : $signed(_GEN_964); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_966 = 7'h2f == data1Frac_7 ? $signed(8'sh32) : $signed(_GEN_965); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_967 = 7'h30 == data1Frac_7 ? $signed(8'sh31) : $signed(_GEN_966); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_968 = 7'h31 == data1Frac_7 ? $signed(8'sh31) : $signed(_GEN_967); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_969 = 7'h32 == data1Frac_7 ? $signed(8'sh31) : $signed(_GEN_968); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_970 = 7'h33 == data1Frac_7 ? $signed(8'sh31) : $signed(_GEN_969); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_971 = 7'h34 == data1Frac_7 ? $signed(8'sh30) : $signed(_GEN_970); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_972 = 7'h35 == data1Frac_7 ? $signed(8'sh30) : $signed(_GEN_971); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_973 = 7'h36 == data1Frac_7 ? $signed(8'sh30) : $signed(_GEN_972); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_974 = 7'h37 == data1Frac_7 ? $signed(8'sh30) : $signed(_GEN_973); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_975 = 7'h38 == data1Frac_7 ? $signed(8'sh2f) : $signed(_GEN_974); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_976 = 7'h39 == data1Frac_7 ? $signed(8'sh2f) : $signed(_GEN_975); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_977 = 7'h3a == data1Frac_7 ? $signed(8'sh2f) : $signed(_GEN_976); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_978 = 7'h3b == data1Frac_7 ? $signed(8'sh2e) : $signed(_GEN_977); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_979 = 7'h3c == data1Frac_7 ? $signed(8'sh2e) : $signed(_GEN_978); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_980 = 7'h3d == data1Frac_7 ? $signed(8'sh2e) : $signed(_GEN_979); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_981 = 7'h3e == data1Frac_7 ? $signed(8'sh2e) : $signed(_GEN_980); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_982 = 7'h3f == data1Frac_7 ? $signed(8'sh2e) : $signed(_GEN_981); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_983 = 7'h40 == data1Frac_7 ? $signed(8'sh2d) : $signed(_GEN_982); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_984 = 7'h41 == data1Frac_7 ? $signed(8'sh2d) : $signed(_GEN_983); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_985 = 7'h42 == data1Frac_7 ? $signed(8'sh2d) : $signed(_GEN_984); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_986 = 7'h43 == data1Frac_7 ? $signed(8'sh2d) : $signed(_GEN_985); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_987 = 7'h44 == data1Frac_7 ? $signed(8'sh2c) : $signed(_GEN_986); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_988 = 7'h45 == data1Frac_7 ? $signed(8'sh2c) : $signed(_GEN_987); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_989 = 7'h46 == data1Frac_7 ? $signed(8'sh2c) : $signed(_GEN_988); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_990 = 7'h47 == data1Frac_7 ? $signed(8'sh2c) : $signed(_GEN_989); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_991 = 7'h48 == data1Frac_7 ? $signed(8'sh2b) : $signed(_GEN_990); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_992 = 7'h49 == data1Frac_7 ? $signed(8'sh2b) : $signed(_GEN_991); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_993 = 7'h4a == data1Frac_7 ? $signed(8'sh2b) : $signed(_GEN_992); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_994 = 7'h4b == data1Frac_7 ? $signed(8'sh2b) : $signed(_GEN_993); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_995 = 7'h4c == data1Frac_7 ? $signed(8'sh2a) : $signed(_GEN_994); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_996 = 7'h4d == data1Frac_7 ? $signed(8'sh2a) : $signed(_GEN_995); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_997 = 7'h4e == data1Frac_7 ? $signed(8'sh2a) : $signed(_GEN_996); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_998 = 7'h4f == data1Frac_7 ? $signed(8'sh2a) : $signed(_GEN_997); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_999 = 7'h50 == data1Frac_7 ? $signed(8'sh29) : $signed(_GEN_998); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1000 = 7'h51 == data1Frac_7 ? $signed(8'sh29) : $signed(_GEN_999); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1001 = 7'h52 == data1Frac_7 ? $signed(8'sh29) : $signed(_GEN_1000); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1002 = 7'h53 == data1Frac_7 ? $signed(8'sh29) : $signed(_GEN_1001); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1003 = 7'h54 == data1Frac_7 ? $signed(8'sh29) : $signed(_GEN_1002); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1004 = 7'h55 == data1Frac_7 ? $signed(8'sh28) : $signed(_GEN_1003); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1005 = 7'h56 == data1Frac_7 ? $signed(8'sh28) : $signed(_GEN_1004); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1006 = 7'h57 == data1Frac_7 ? $signed(8'sh28) : $signed(_GEN_1005); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1007 = 7'h58 == data1Frac_7 ? $signed(8'sh28) : $signed(_GEN_1006); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1008 = 7'h59 == data1Frac_7 ? $signed(8'sh28) : $signed(_GEN_1007); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1009 = 7'h5a == data1Frac_7 ? $signed(8'sh27) : $signed(_GEN_1008); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1010 = 7'h5b == data1Frac_7 ? $signed(8'sh27) : $signed(_GEN_1009); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1011 = 7'h5c == data1Frac_7 ? $signed(8'sh27) : $signed(_GEN_1010); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1012 = 7'h5d == data1Frac_7 ? $signed(8'sh27) : $signed(_GEN_1011); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1013 = 7'h5e == data1Frac_7 ? $signed(8'sh26) : $signed(_GEN_1012); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1014 = 7'h5f == data1Frac_7 ? $signed(8'sh26) : $signed(_GEN_1013); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1015 = 7'h60 == data1Frac_7 ? $signed(8'sh26) : $signed(_GEN_1014); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1016 = 7'h61 == data1Frac_7 ? $signed(8'sh26) : $signed(_GEN_1015); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1017 = 7'h62 == data1Frac_7 ? $signed(8'sh26) : $signed(_GEN_1016); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1018 = 7'h63 == data1Frac_7 ? $signed(8'sh25) : $signed(_GEN_1017); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1019 = 7'h64 == data1Frac_7 ? $signed(8'sh25) : $signed(_GEN_1018); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1020 = 7'h65 == data1Frac_7 ? $signed(8'sh25) : $signed(_GEN_1019); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1021 = 7'h66 == data1Frac_7 ? $signed(8'sh25) : $signed(_GEN_1020); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1022 = 7'h67 == data1Frac_7 ? $signed(8'sh25) : $signed(_GEN_1021); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1023 = 7'h68 == data1Frac_7 ? $signed(8'sh24) : $signed(_GEN_1022); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1024 = 7'h69 == data1Frac_7 ? $signed(8'sh24) : $signed(_GEN_1023); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1025 = 7'h6a == data1Frac_7 ? $signed(8'sh24) : $signed(_GEN_1024); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1026 = 7'h6b == data1Frac_7 ? $signed(8'sh24) : $signed(_GEN_1025); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1027 = 7'h6c == data1Frac_7 ? $signed(8'sh24) : $signed(_GEN_1026); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1028 = 7'h6d == data1Frac_7 ? $signed(8'sh23) : $signed(_GEN_1027); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1029 = 7'h6e == data1Frac_7 ? $signed(8'sh23) : $signed(_GEN_1028); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1030 = 7'h6f == data1Frac_7 ? $signed(8'sh23) : $signed(_GEN_1029); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1031 = 7'h70 == data1Frac_7 ? $signed(8'sh23) : $signed(_GEN_1030); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1032 = 7'h71 == data1Frac_7 ? $signed(8'sh23) : $signed(_GEN_1031); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1033 = 7'h72 == data1Frac_7 ? $signed(8'sh23) : $signed(_GEN_1032); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1034 = 7'h73 == data1Frac_7 ? $signed(8'sh22) : $signed(_GEN_1033); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1035 = 7'h74 == data1Frac_7 ? $signed(8'sh22) : $signed(_GEN_1034); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1036 = 7'h75 == data1Frac_7 ? $signed(8'sh22) : $signed(_GEN_1035); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1037 = 7'h76 == data1Frac_7 ? $signed(8'sh22) : $signed(_GEN_1036); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1038 = 7'h77 == data1Frac_7 ? $signed(8'sh22) : $signed(_GEN_1037); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1039 = 7'h78 == data1Frac_7 ? $signed(8'sh21) : $signed(_GEN_1038); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1040 = 7'h79 == data1Frac_7 ? $signed(8'sh21) : $signed(_GEN_1039); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1041 = 7'h7a == data1Frac_7 ? $signed(8'sh21) : $signed(_GEN_1040); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1042 = 7'h7b == data1Frac_7 ? $signed(8'sh21) : $signed(_GEN_1041); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1043 = 7'h7c == data1Frac_7 ? $signed(8'sh21) : $signed(_GEN_1042); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1044 = 7'h7d == data1Frac_7 ? $signed(8'sh21) : $signed(_GEN_1043); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1045 = 7'h7e == data1Frac_7 ? $signed(8'sh20) : $signed(_GEN_1044); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1046 = 7'h7f == data1Frac_7 ? $signed(8'sh20) : $signed(_GEN_1045); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_23 = $signed(_GEN_1046) >>> data1Int_7; // @[exponent.scala 38:85]
  reg [7:0] data2_7; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1050 = 7'h2 == data1Frac_8 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1051 = 7'h3 == data1Frac_8 ? $signed(8'sh3f) : $signed(_GEN_1050); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1052 = 7'h4 == data1Frac_8 ? $signed(8'sh3f) : $signed(_GEN_1051); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1053 = 7'h5 == data1Frac_8 ? $signed(8'sh3e) : $signed(_GEN_1052); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1054 = 7'h6 == data1Frac_8 ? $signed(8'sh3e) : $signed(_GEN_1053); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1055 = 7'h7 == data1Frac_8 ? $signed(8'sh3e) : $signed(_GEN_1054); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1056 = 7'h8 == data1Frac_8 ? $signed(8'sh3d) : $signed(_GEN_1055); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1057 = 7'h9 == data1Frac_8 ? $signed(8'sh3d) : $signed(_GEN_1056); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1058 = 7'ha == data1Frac_8 ? $signed(8'sh3d) : $signed(_GEN_1057); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1059 = 7'hb == data1Frac_8 ? $signed(8'sh3c) : $signed(_GEN_1058); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1060 = 7'hc == data1Frac_8 ? $signed(8'sh3c) : $signed(_GEN_1059); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1061 = 7'hd == data1Frac_8 ? $signed(8'sh3c) : $signed(_GEN_1060); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1062 = 7'he == data1Frac_8 ? $signed(8'sh3b) : $signed(_GEN_1061); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1063 = 7'hf == data1Frac_8 ? $signed(8'sh3b) : $signed(_GEN_1062); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1064 = 7'h10 == data1Frac_8 ? $signed(8'sh3b) : $signed(_GEN_1063); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1065 = 7'h11 == data1Frac_8 ? $signed(8'sh3a) : $signed(_GEN_1064); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1066 = 7'h12 == data1Frac_8 ? $signed(8'sh3a) : $signed(_GEN_1065); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1067 = 7'h13 == data1Frac_8 ? $signed(8'sh3a) : $signed(_GEN_1066); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1068 = 7'h14 == data1Frac_8 ? $signed(8'sh39) : $signed(_GEN_1067); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1069 = 7'h15 == data1Frac_8 ? $signed(8'sh39) : $signed(_GEN_1068); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1070 = 7'h16 == data1Frac_8 ? $signed(8'sh39) : $signed(_GEN_1069); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1071 = 7'h17 == data1Frac_8 ? $signed(8'sh39) : $signed(_GEN_1070); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1072 = 7'h18 == data1Frac_8 ? $signed(8'sh38) : $signed(_GEN_1071); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1073 = 7'h19 == data1Frac_8 ? $signed(8'sh38) : $signed(_GEN_1072); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1074 = 7'h1a == data1Frac_8 ? $signed(8'sh38) : $signed(_GEN_1073); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1075 = 7'h1b == data1Frac_8 ? $signed(8'sh37) : $signed(_GEN_1074); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1076 = 7'h1c == data1Frac_8 ? $signed(8'sh37) : $signed(_GEN_1075); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1077 = 7'h1d == data1Frac_8 ? $signed(8'sh37) : $signed(_GEN_1076); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1078 = 7'h1e == data1Frac_8 ? $signed(8'sh36) : $signed(_GEN_1077); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1079 = 7'h1f == data1Frac_8 ? $signed(8'sh36) : $signed(_GEN_1078); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1080 = 7'h20 == data1Frac_8 ? $signed(8'sh36) : $signed(_GEN_1079); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1081 = 7'h21 == data1Frac_8 ? $signed(8'sh36) : $signed(_GEN_1080); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1082 = 7'h22 == data1Frac_8 ? $signed(8'sh35) : $signed(_GEN_1081); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1083 = 7'h23 == data1Frac_8 ? $signed(8'sh35) : $signed(_GEN_1082); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1084 = 7'h24 == data1Frac_8 ? $signed(8'sh35) : $signed(_GEN_1083); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1085 = 7'h25 == data1Frac_8 ? $signed(8'sh34) : $signed(_GEN_1084); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1086 = 7'h26 == data1Frac_8 ? $signed(8'sh34) : $signed(_GEN_1085); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1087 = 7'h27 == data1Frac_8 ? $signed(8'sh34) : $signed(_GEN_1086); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1088 = 7'h28 == data1Frac_8 ? $signed(8'sh34) : $signed(_GEN_1087); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1089 = 7'h29 == data1Frac_8 ? $signed(8'sh33) : $signed(_GEN_1088); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1090 = 7'h2a == data1Frac_8 ? $signed(8'sh33) : $signed(_GEN_1089); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1091 = 7'h2b == data1Frac_8 ? $signed(8'sh33) : $signed(_GEN_1090); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1092 = 7'h2c == data1Frac_8 ? $signed(8'sh32) : $signed(_GEN_1091); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1093 = 7'h2d == data1Frac_8 ? $signed(8'sh32) : $signed(_GEN_1092); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1094 = 7'h2e == data1Frac_8 ? $signed(8'sh32) : $signed(_GEN_1093); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1095 = 7'h2f == data1Frac_8 ? $signed(8'sh32) : $signed(_GEN_1094); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1096 = 7'h30 == data1Frac_8 ? $signed(8'sh31) : $signed(_GEN_1095); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1097 = 7'h31 == data1Frac_8 ? $signed(8'sh31) : $signed(_GEN_1096); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1098 = 7'h32 == data1Frac_8 ? $signed(8'sh31) : $signed(_GEN_1097); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1099 = 7'h33 == data1Frac_8 ? $signed(8'sh31) : $signed(_GEN_1098); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1100 = 7'h34 == data1Frac_8 ? $signed(8'sh30) : $signed(_GEN_1099); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1101 = 7'h35 == data1Frac_8 ? $signed(8'sh30) : $signed(_GEN_1100); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1102 = 7'h36 == data1Frac_8 ? $signed(8'sh30) : $signed(_GEN_1101); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1103 = 7'h37 == data1Frac_8 ? $signed(8'sh30) : $signed(_GEN_1102); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1104 = 7'h38 == data1Frac_8 ? $signed(8'sh2f) : $signed(_GEN_1103); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1105 = 7'h39 == data1Frac_8 ? $signed(8'sh2f) : $signed(_GEN_1104); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1106 = 7'h3a == data1Frac_8 ? $signed(8'sh2f) : $signed(_GEN_1105); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1107 = 7'h3b == data1Frac_8 ? $signed(8'sh2e) : $signed(_GEN_1106); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1108 = 7'h3c == data1Frac_8 ? $signed(8'sh2e) : $signed(_GEN_1107); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1109 = 7'h3d == data1Frac_8 ? $signed(8'sh2e) : $signed(_GEN_1108); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1110 = 7'h3e == data1Frac_8 ? $signed(8'sh2e) : $signed(_GEN_1109); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1111 = 7'h3f == data1Frac_8 ? $signed(8'sh2e) : $signed(_GEN_1110); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1112 = 7'h40 == data1Frac_8 ? $signed(8'sh2d) : $signed(_GEN_1111); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1113 = 7'h41 == data1Frac_8 ? $signed(8'sh2d) : $signed(_GEN_1112); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1114 = 7'h42 == data1Frac_8 ? $signed(8'sh2d) : $signed(_GEN_1113); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1115 = 7'h43 == data1Frac_8 ? $signed(8'sh2d) : $signed(_GEN_1114); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1116 = 7'h44 == data1Frac_8 ? $signed(8'sh2c) : $signed(_GEN_1115); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1117 = 7'h45 == data1Frac_8 ? $signed(8'sh2c) : $signed(_GEN_1116); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1118 = 7'h46 == data1Frac_8 ? $signed(8'sh2c) : $signed(_GEN_1117); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1119 = 7'h47 == data1Frac_8 ? $signed(8'sh2c) : $signed(_GEN_1118); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1120 = 7'h48 == data1Frac_8 ? $signed(8'sh2b) : $signed(_GEN_1119); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1121 = 7'h49 == data1Frac_8 ? $signed(8'sh2b) : $signed(_GEN_1120); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1122 = 7'h4a == data1Frac_8 ? $signed(8'sh2b) : $signed(_GEN_1121); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1123 = 7'h4b == data1Frac_8 ? $signed(8'sh2b) : $signed(_GEN_1122); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1124 = 7'h4c == data1Frac_8 ? $signed(8'sh2a) : $signed(_GEN_1123); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1125 = 7'h4d == data1Frac_8 ? $signed(8'sh2a) : $signed(_GEN_1124); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1126 = 7'h4e == data1Frac_8 ? $signed(8'sh2a) : $signed(_GEN_1125); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1127 = 7'h4f == data1Frac_8 ? $signed(8'sh2a) : $signed(_GEN_1126); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1128 = 7'h50 == data1Frac_8 ? $signed(8'sh29) : $signed(_GEN_1127); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1129 = 7'h51 == data1Frac_8 ? $signed(8'sh29) : $signed(_GEN_1128); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1130 = 7'h52 == data1Frac_8 ? $signed(8'sh29) : $signed(_GEN_1129); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1131 = 7'h53 == data1Frac_8 ? $signed(8'sh29) : $signed(_GEN_1130); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1132 = 7'h54 == data1Frac_8 ? $signed(8'sh29) : $signed(_GEN_1131); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1133 = 7'h55 == data1Frac_8 ? $signed(8'sh28) : $signed(_GEN_1132); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1134 = 7'h56 == data1Frac_8 ? $signed(8'sh28) : $signed(_GEN_1133); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1135 = 7'h57 == data1Frac_8 ? $signed(8'sh28) : $signed(_GEN_1134); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1136 = 7'h58 == data1Frac_8 ? $signed(8'sh28) : $signed(_GEN_1135); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1137 = 7'h59 == data1Frac_8 ? $signed(8'sh28) : $signed(_GEN_1136); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1138 = 7'h5a == data1Frac_8 ? $signed(8'sh27) : $signed(_GEN_1137); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1139 = 7'h5b == data1Frac_8 ? $signed(8'sh27) : $signed(_GEN_1138); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1140 = 7'h5c == data1Frac_8 ? $signed(8'sh27) : $signed(_GEN_1139); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1141 = 7'h5d == data1Frac_8 ? $signed(8'sh27) : $signed(_GEN_1140); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1142 = 7'h5e == data1Frac_8 ? $signed(8'sh26) : $signed(_GEN_1141); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1143 = 7'h5f == data1Frac_8 ? $signed(8'sh26) : $signed(_GEN_1142); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1144 = 7'h60 == data1Frac_8 ? $signed(8'sh26) : $signed(_GEN_1143); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1145 = 7'h61 == data1Frac_8 ? $signed(8'sh26) : $signed(_GEN_1144); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1146 = 7'h62 == data1Frac_8 ? $signed(8'sh26) : $signed(_GEN_1145); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1147 = 7'h63 == data1Frac_8 ? $signed(8'sh25) : $signed(_GEN_1146); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1148 = 7'h64 == data1Frac_8 ? $signed(8'sh25) : $signed(_GEN_1147); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1149 = 7'h65 == data1Frac_8 ? $signed(8'sh25) : $signed(_GEN_1148); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1150 = 7'h66 == data1Frac_8 ? $signed(8'sh25) : $signed(_GEN_1149); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1151 = 7'h67 == data1Frac_8 ? $signed(8'sh25) : $signed(_GEN_1150); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1152 = 7'h68 == data1Frac_8 ? $signed(8'sh24) : $signed(_GEN_1151); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1153 = 7'h69 == data1Frac_8 ? $signed(8'sh24) : $signed(_GEN_1152); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1154 = 7'h6a == data1Frac_8 ? $signed(8'sh24) : $signed(_GEN_1153); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1155 = 7'h6b == data1Frac_8 ? $signed(8'sh24) : $signed(_GEN_1154); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1156 = 7'h6c == data1Frac_8 ? $signed(8'sh24) : $signed(_GEN_1155); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1157 = 7'h6d == data1Frac_8 ? $signed(8'sh23) : $signed(_GEN_1156); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1158 = 7'h6e == data1Frac_8 ? $signed(8'sh23) : $signed(_GEN_1157); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1159 = 7'h6f == data1Frac_8 ? $signed(8'sh23) : $signed(_GEN_1158); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1160 = 7'h70 == data1Frac_8 ? $signed(8'sh23) : $signed(_GEN_1159); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1161 = 7'h71 == data1Frac_8 ? $signed(8'sh23) : $signed(_GEN_1160); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1162 = 7'h72 == data1Frac_8 ? $signed(8'sh23) : $signed(_GEN_1161); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1163 = 7'h73 == data1Frac_8 ? $signed(8'sh22) : $signed(_GEN_1162); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1164 = 7'h74 == data1Frac_8 ? $signed(8'sh22) : $signed(_GEN_1163); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1165 = 7'h75 == data1Frac_8 ? $signed(8'sh22) : $signed(_GEN_1164); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1166 = 7'h76 == data1Frac_8 ? $signed(8'sh22) : $signed(_GEN_1165); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1167 = 7'h77 == data1Frac_8 ? $signed(8'sh22) : $signed(_GEN_1166); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1168 = 7'h78 == data1Frac_8 ? $signed(8'sh21) : $signed(_GEN_1167); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1169 = 7'h79 == data1Frac_8 ? $signed(8'sh21) : $signed(_GEN_1168); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1170 = 7'h7a == data1Frac_8 ? $signed(8'sh21) : $signed(_GEN_1169); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1171 = 7'h7b == data1Frac_8 ? $signed(8'sh21) : $signed(_GEN_1170); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1172 = 7'h7c == data1Frac_8 ? $signed(8'sh21) : $signed(_GEN_1171); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1173 = 7'h7d == data1Frac_8 ? $signed(8'sh21) : $signed(_GEN_1172); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1174 = 7'h7e == data1Frac_8 ? $signed(8'sh20) : $signed(_GEN_1173); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1175 = 7'h7f == data1Frac_8 ? $signed(8'sh20) : $signed(_GEN_1174); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_26 = $signed(_GEN_1175) >>> data1Int_8; // @[exponent.scala 38:85]
  reg [7:0] data2_8; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1179 = 7'h2 == data1Frac_9 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1180 = 7'h3 == data1Frac_9 ? $signed(8'sh3f) : $signed(_GEN_1179); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1181 = 7'h4 == data1Frac_9 ? $signed(8'sh3f) : $signed(_GEN_1180); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1182 = 7'h5 == data1Frac_9 ? $signed(8'sh3e) : $signed(_GEN_1181); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1183 = 7'h6 == data1Frac_9 ? $signed(8'sh3e) : $signed(_GEN_1182); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1184 = 7'h7 == data1Frac_9 ? $signed(8'sh3e) : $signed(_GEN_1183); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1185 = 7'h8 == data1Frac_9 ? $signed(8'sh3d) : $signed(_GEN_1184); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1186 = 7'h9 == data1Frac_9 ? $signed(8'sh3d) : $signed(_GEN_1185); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1187 = 7'ha == data1Frac_9 ? $signed(8'sh3d) : $signed(_GEN_1186); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1188 = 7'hb == data1Frac_9 ? $signed(8'sh3c) : $signed(_GEN_1187); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1189 = 7'hc == data1Frac_9 ? $signed(8'sh3c) : $signed(_GEN_1188); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1190 = 7'hd == data1Frac_9 ? $signed(8'sh3c) : $signed(_GEN_1189); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1191 = 7'he == data1Frac_9 ? $signed(8'sh3b) : $signed(_GEN_1190); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1192 = 7'hf == data1Frac_9 ? $signed(8'sh3b) : $signed(_GEN_1191); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1193 = 7'h10 == data1Frac_9 ? $signed(8'sh3b) : $signed(_GEN_1192); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1194 = 7'h11 == data1Frac_9 ? $signed(8'sh3a) : $signed(_GEN_1193); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1195 = 7'h12 == data1Frac_9 ? $signed(8'sh3a) : $signed(_GEN_1194); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1196 = 7'h13 == data1Frac_9 ? $signed(8'sh3a) : $signed(_GEN_1195); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1197 = 7'h14 == data1Frac_9 ? $signed(8'sh39) : $signed(_GEN_1196); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1198 = 7'h15 == data1Frac_9 ? $signed(8'sh39) : $signed(_GEN_1197); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1199 = 7'h16 == data1Frac_9 ? $signed(8'sh39) : $signed(_GEN_1198); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1200 = 7'h17 == data1Frac_9 ? $signed(8'sh39) : $signed(_GEN_1199); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1201 = 7'h18 == data1Frac_9 ? $signed(8'sh38) : $signed(_GEN_1200); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1202 = 7'h19 == data1Frac_9 ? $signed(8'sh38) : $signed(_GEN_1201); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1203 = 7'h1a == data1Frac_9 ? $signed(8'sh38) : $signed(_GEN_1202); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1204 = 7'h1b == data1Frac_9 ? $signed(8'sh37) : $signed(_GEN_1203); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1205 = 7'h1c == data1Frac_9 ? $signed(8'sh37) : $signed(_GEN_1204); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1206 = 7'h1d == data1Frac_9 ? $signed(8'sh37) : $signed(_GEN_1205); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1207 = 7'h1e == data1Frac_9 ? $signed(8'sh36) : $signed(_GEN_1206); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1208 = 7'h1f == data1Frac_9 ? $signed(8'sh36) : $signed(_GEN_1207); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1209 = 7'h20 == data1Frac_9 ? $signed(8'sh36) : $signed(_GEN_1208); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1210 = 7'h21 == data1Frac_9 ? $signed(8'sh36) : $signed(_GEN_1209); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1211 = 7'h22 == data1Frac_9 ? $signed(8'sh35) : $signed(_GEN_1210); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1212 = 7'h23 == data1Frac_9 ? $signed(8'sh35) : $signed(_GEN_1211); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1213 = 7'h24 == data1Frac_9 ? $signed(8'sh35) : $signed(_GEN_1212); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1214 = 7'h25 == data1Frac_9 ? $signed(8'sh34) : $signed(_GEN_1213); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1215 = 7'h26 == data1Frac_9 ? $signed(8'sh34) : $signed(_GEN_1214); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1216 = 7'h27 == data1Frac_9 ? $signed(8'sh34) : $signed(_GEN_1215); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1217 = 7'h28 == data1Frac_9 ? $signed(8'sh34) : $signed(_GEN_1216); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1218 = 7'h29 == data1Frac_9 ? $signed(8'sh33) : $signed(_GEN_1217); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1219 = 7'h2a == data1Frac_9 ? $signed(8'sh33) : $signed(_GEN_1218); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1220 = 7'h2b == data1Frac_9 ? $signed(8'sh33) : $signed(_GEN_1219); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1221 = 7'h2c == data1Frac_9 ? $signed(8'sh32) : $signed(_GEN_1220); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1222 = 7'h2d == data1Frac_9 ? $signed(8'sh32) : $signed(_GEN_1221); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1223 = 7'h2e == data1Frac_9 ? $signed(8'sh32) : $signed(_GEN_1222); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1224 = 7'h2f == data1Frac_9 ? $signed(8'sh32) : $signed(_GEN_1223); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1225 = 7'h30 == data1Frac_9 ? $signed(8'sh31) : $signed(_GEN_1224); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1226 = 7'h31 == data1Frac_9 ? $signed(8'sh31) : $signed(_GEN_1225); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1227 = 7'h32 == data1Frac_9 ? $signed(8'sh31) : $signed(_GEN_1226); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1228 = 7'h33 == data1Frac_9 ? $signed(8'sh31) : $signed(_GEN_1227); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1229 = 7'h34 == data1Frac_9 ? $signed(8'sh30) : $signed(_GEN_1228); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1230 = 7'h35 == data1Frac_9 ? $signed(8'sh30) : $signed(_GEN_1229); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1231 = 7'h36 == data1Frac_9 ? $signed(8'sh30) : $signed(_GEN_1230); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1232 = 7'h37 == data1Frac_9 ? $signed(8'sh30) : $signed(_GEN_1231); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1233 = 7'h38 == data1Frac_9 ? $signed(8'sh2f) : $signed(_GEN_1232); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1234 = 7'h39 == data1Frac_9 ? $signed(8'sh2f) : $signed(_GEN_1233); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1235 = 7'h3a == data1Frac_9 ? $signed(8'sh2f) : $signed(_GEN_1234); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1236 = 7'h3b == data1Frac_9 ? $signed(8'sh2e) : $signed(_GEN_1235); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1237 = 7'h3c == data1Frac_9 ? $signed(8'sh2e) : $signed(_GEN_1236); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1238 = 7'h3d == data1Frac_9 ? $signed(8'sh2e) : $signed(_GEN_1237); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1239 = 7'h3e == data1Frac_9 ? $signed(8'sh2e) : $signed(_GEN_1238); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1240 = 7'h3f == data1Frac_9 ? $signed(8'sh2e) : $signed(_GEN_1239); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1241 = 7'h40 == data1Frac_9 ? $signed(8'sh2d) : $signed(_GEN_1240); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1242 = 7'h41 == data1Frac_9 ? $signed(8'sh2d) : $signed(_GEN_1241); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1243 = 7'h42 == data1Frac_9 ? $signed(8'sh2d) : $signed(_GEN_1242); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1244 = 7'h43 == data1Frac_9 ? $signed(8'sh2d) : $signed(_GEN_1243); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1245 = 7'h44 == data1Frac_9 ? $signed(8'sh2c) : $signed(_GEN_1244); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1246 = 7'h45 == data1Frac_9 ? $signed(8'sh2c) : $signed(_GEN_1245); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1247 = 7'h46 == data1Frac_9 ? $signed(8'sh2c) : $signed(_GEN_1246); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1248 = 7'h47 == data1Frac_9 ? $signed(8'sh2c) : $signed(_GEN_1247); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1249 = 7'h48 == data1Frac_9 ? $signed(8'sh2b) : $signed(_GEN_1248); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1250 = 7'h49 == data1Frac_9 ? $signed(8'sh2b) : $signed(_GEN_1249); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1251 = 7'h4a == data1Frac_9 ? $signed(8'sh2b) : $signed(_GEN_1250); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1252 = 7'h4b == data1Frac_9 ? $signed(8'sh2b) : $signed(_GEN_1251); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1253 = 7'h4c == data1Frac_9 ? $signed(8'sh2a) : $signed(_GEN_1252); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1254 = 7'h4d == data1Frac_9 ? $signed(8'sh2a) : $signed(_GEN_1253); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1255 = 7'h4e == data1Frac_9 ? $signed(8'sh2a) : $signed(_GEN_1254); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1256 = 7'h4f == data1Frac_9 ? $signed(8'sh2a) : $signed(_GEN_1255); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1257 = 7'h50 == data1Frac_9 ? $signed(8'sh29) : $signed(_GEN_1256); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1258 = 7'h51 == data1Frac_9 ? $signed(8'sh29) : $signed(_GEN_1257); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1259 = 7'h52 == data1Frac_9 ? $signed(8'sh29) : $signed(_GEN_1258); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1260 = 7'h53 == data1Frac_9 ? $signed(8'sh29) : $signed(_GEN_1259); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1261 = 7'h54 == data1Frac_9 ? $signed(8'sh29) : $signed(_GEN_1260); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1262 = 7'h55 == data1Frac_9 ? $signed(8'sh28) : $signed(_GEN_1261); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1263 = 7'h56 == data1Frac_9 ? $signed(8'sh28) : $signed(_GEN_1262); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1264 = 7'h57 == data1Frac_9 ? $signed(8'sh28) : $signed(_GEN_1263); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1265 = 7'h58 == data1Frac_9 ? $signed(8'sh28) : $signed(_GEN_1264); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1266 = 7'h59 == data1Frac_9 ? $signed(8'sh28) : $signed(_GEN_1265); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1267 = 7'h5a == data1Frac_9 ? $signed(8'sh27) : $signed(_GEN_1266); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1268 = 7'h5b == data1Frac_9 ? $signed(8'sh27) : $signed(_GEN_1267); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1269 = 7'h5c == data1Frac_9 ? $signed(8'sh27) : $signed(_GEN_1268); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1270 = 7'h5d == data1Frac_9 ? $signed(8'sh27) : $signed(_GEN_1269); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1271 = 7'h5e == data1Frac_9 ? $signed(8'sh26) : $signed(_GEN_1270); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1272 = 7'h5f == data1Frac_9 ? $signed(8'sh26) : $signed(_GEN_1271); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1273 = 7'h60 == data1Frac_9 ? $signed(8'sh26) : $signed(_GEN_1272); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1274 = 7'h61 == data1Frac_9 ? $signed(8'sh26) : $signed(_GEN_1273); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1275 = 7'h62 == data1Frac_9 ? $signed(8'sh26) : $signed(_GEN_1274); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1276 = 7'h63 == data1Frac_9 ? $signed(8'sh25) : $signed(_GEN_1275); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1277 = 7'h64 == data1Frac_9 ? $signed(8'sh25) : $signed(_GEN_1276); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1278 = 7'h65 == data1Frac_9 ? $signed(8'sh25) : $signed(_GEN_1277); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1279 = 7'h66 == data1Frac_9 ? $signed(8'sh25) : $signed(_GEN_1278); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1280 = 7'h67 == data1Frac_9 ? $signed(8'sh25) : $signed(_GEN_1279); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1281 = 7'h68 == data1Frac_9 ? $signed(8'sh24) : $signed(_GEN_1280); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1282 = 7'h69 == data1Frac_9 ? $signed(8'sh24) : $signed(_GEN_1281); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1283 = 7'h6a == data1Frac_9 ? $signed(8'sh24) : $signed(_GEN_1282); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1284 = 7'h6b == data1Frac_9 ? $signed(8'sh24) : $signed(_GEN_1283); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1285 = 7'h6c == data1Frac_9 ? $signed(8'sh24) : $signed(_GEN_1284); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1286 = 7'h6d == data1Frac_9 ? $signed(8'sh23) : $signed(_GEN_1285); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1287 = 7'h6e == data1Frac_9 ? $signed(8'sh23) : $signed(_GEN_1286); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1288 = 7'h6f == data1Frac_9 ? $signed(8'sh23) : $signed(_GEN_1287); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1289 = 7'h70 == data1Frac_9 ? $signed(8'sh23) : $signed(_GEN_1288); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1290 = 7'h71 == data1Frac_9 ? $signed(8'sh23) : $signed(_GEN_1289); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1291 = 7'h72 == data1Frac_9 ? $signed(8'sh23) : $signed(_GEN_1290); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1292 = 7'h73 == data1Frac_9 ? $signed(8'sh22) : $signed(_GEN_1291); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1293 = 7'h74 == data1Frac_9 ? $signed(8'sh22) : $signed(_GEN_1292); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1294 = 7'h75 == data1Frac_9 ? $signed(8'sh22) : $signed(_GEN_1293); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1295 = 7'h76 == data1Frac_9 ? $signed(8'sh22) : $signed(_GEN_1294); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1296 = 7'h77 == data1Frac_9 ? $signed(8'sh22) : $signed(_GEN_1295); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1297 = 7'h78 == data1Frac_9 ? $signed(8'sh21) : $signed(_GEN_1296); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1298 = 7'h79 == data1Frac_9 ? $signed(8'sh21) : $signed(_GEN_1297); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1299 = 7'h7a == data1Frac_9 ? $signed(8'sh21) : $signed(_GEN_1298); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1300 = 7'h7b == data1Frac_9 ? $signed(8'sh21) : $signed(_GEN_1299); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1301 = 7'h7c == data1Frac_9 ? $signed(8'sh21) : $signed(_GEN_1300); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1302 = 7'h7d == data1Frac_9 ? $signed(8'sh21) : $signed(_GEN_1301); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1303 = 7'h7e == data1Frac_9 ? $signed(8'sh20) : $signed(_GEN_1302); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1304 = 7'h7f == data1Frac_9 ? $signed(8'sh20) : $signed(_GEN_1303); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_29 = $signed(_GEN_1304) >>> data1Int_9; // @[exponent.scala 38:85]
  reg [7:0] data2_9; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1308 = 7'h2 == data1Frac_10 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1309 = 7'h3 == data1Frac_10 ? $signed(8'sh3f) : $signed(_GEN_1308); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1310 = 7'h4 == data1Frac_10 ? $signed(8'sh3f) : $signed(_GEN_1309); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1311 = 7'h5 == data1Frac_10 ? $signed(8'sh3e) : $signed(_GEN_1310); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1312 = 7'h6 == data1Frac_10 ? $signed(8'sh3e) : $signed(_GEN_1311); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1313 = 7'h7 == data1Frac_10 ? $signed(8'sh3e) : $signed(_GEN_1312); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1314 = 7'h8 == data1Frac_10 ? $signed(8'sh3d) : $signed(_GEN_1313); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1315 = 7'h9 == data1Frac_10 ? $signed(8'sh3d) : $signed(_GEN_1314); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1316 = 7'ha == data1Frac_10 ? $signed(8'sh3d) : $signed(_GEN_1315); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1317 = 7'hb == data1Frac_10 ? $signed(8'sh3c) : $signed(_GEN_1316); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1318 = 7'hc == data1Frac_10 ? $signed(8'sh3c) : $signed(_GEN_1317); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1319 = 7'hd == data1Frac_10 ? $signed(8'sh3c) : $signed(_GEN_1318); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1320 = 7'he == data1Frac_10 ? $signed(8'sh3b) : $signed(_GEN_1319); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1321 = 7'hf == data1Frac_10 ? $signed(8'sh3b) : $signed(_GEN_1320); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1322 = 7'h10 == data1Frac_10 ? $signed(8'sh3b) : $signed(_GEN_1321); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1323 = 7'h11 == data1Frac_10 ? $signed(8'sh3a) : $signed(_GEN_1322); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1324 = 7'h12 == data1Frac_10 ? $signed(8'sh3a) : $signed(_GEN_1323); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1325 = 7'h13 == data1Frac_10 ? $signed(8'sh3a) : $signed(_GEN_1324); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1326 = 7'h14 == data1Frac_10 ? $signed(8'sh39) : $signed(_GEN_1325); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1327 = 7'h15 == data1Frac_10 ? $signed(8'sh39) : $signed(_GEN_1326); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1328 = 7'h16 == data1Frac_10 ? $signed(8'sh39) : $signed(_GEN_1327); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1329 = 7'h17 == data1Frac_10 ? $signed(8'sh39) : $signed(_GEN_1328); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1330 = 7'h18 == data1Frac_10 ? $signed(8'sh38) : $signed(_GEN_1329); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1331 = 7'h19 == data1Frac_10 ? $signed(8'sh38) : $signed(_GEN_1330); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1332 = 7'h1a == data1Frac_10 ? $signed(8'sh38) : $signed(_GEN_1331); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1333 = 7'h1b == data1Frac_10 ? $signed(8'sh37) : $signed(_GEN_1332); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1334 = 7'h1c == data1Frac_10 ? $signed(8'sh37) : $signed(_GEN_1333); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1335 = 7'h1d == data1Frac_10 ? $signed(8'sh37) : $signed(_GEN_1334); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1336 = 7'h1e == data1Frac_10 ? $signed(8'sh36) : $signed(_GEN_1335); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1337 = 7'h1f == data1Frac_10 ? $signed(8'sh36) : $signed(_GEN_1336); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1338 = 7'h20 == data1Frac_10 ? $signed(8'sh36) : $signed(_GEN_1337); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1339 = 7'h21 == data1Frac_10 ? $signed(8'sh36) : $signed(_GEN_1338); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1340 = 7'h22 == data1Frac_10 ? $signed(8'sh35) : $signed(_GEN_1339); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1341 = 7'h23 == data1Frac_10 ? $signed(8'sh35) : $signed(_GEN_1340); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1342 = 7'h24 == data1Frac_10 ? $signed(8'sh35) : $signed(_GEN_1341); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1343 = 7'h25 == data1Frac_10 ? $signed(8'sh34) : $signed(_GEN_1342); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1344 = 7'h26 == data1Frac_10 ? $signed(8'sh34) : $signed(_GEN_1343); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1345 = 7'h27 == data1Frac_10 ? $signed(8'sh34) : $signed(_GEN_1344); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1346 = 7'h28 == data1Frac_10 ? $signed(8'sh34) : $signed(_GEN_1345); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1347 = 7'h29 == data1Frac_10 ? $signed(8'sh33) : $signed(_GEN_1346); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1348 = 7'h2a == data1Frac_10 ? $signed(8'sh33) : $signed(_GEN_1347); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1349 = 7'h2b == data1Frac_10 ? $signed(8'sh33) : $signed(_GEN_1348); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1350 = 7'h2c == data1Frac_10 ? $signed(8'sh32) : $signed(_GEN_1349); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1351 = 7'h2d == data1Frac_10 ? $signed(8'sh32) : $signed(_GEN_1350); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1352 = 7'h2e == data1Frac_10 ? $signed(8'sh32) : $signed(_GEN_1351); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1353 = 7'h2f == data1Frac_10 ? $signed(8'sh32) : $signed(_GEN_1352); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1354 = 7'h30 == data1Frac_10 ? $signed(8'sh31) : $signed(_GEN_1353); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1355 = 7'h31 == data1Frac_10 ? $signed(8'sh31) : $signed(_GEN_1354); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1356 = 7'h32 == data1Frac_10 ? $signed(8'sh31) : $signed(_GEN_1355); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1357 = 7'h33 == data1Frac_10 ? $signed(8'sh31) : $signed(_GEN_1356); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1358 = 7'h34 == data1Frac_10 ? $signed(8'sh30) : $signed(_GEN_1357); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1359 = 7'h35 == data1Frac_10 ? $signed(8'sh30) : $signed(_GEN_1358); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1360 = 7'h36 == data1Frac_10 ? $signed(8'sh30) : $signed(_GEN_1359); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1361 = 7'h37 == data1Frac_10 ? $signed(8'sh30) : $signed(_GEN_1360); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1362 = 7'h38 == data1Frac_10 ? $signed(8'sh2f) : $signed(_GEN_1361); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1363 = 7'h39 == data1Frac_10 ? $signed(8'sh2f) : $signed(_GEN_1362); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1364 = 7'h3a == data1Frac_10 ? $signed(8'sh2f) : $signed(_GEN_1363); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1365 = 7'h3b == data1Frac_10 ? $signed(8'sh2e) : $signed(_GEN_1364); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1366 = 7'h3c == data1Frac_10 ? $signed(8'sh2e) : $signed(_GEN_1365); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1367 = 7'h3d == data1Frac_10 ? $signed(8'sh2e) : $signed(_GEN_1366); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1368 = 7'h3e == data1Frac_10 ? $signed(8'sh2e) : $signed(_GEN_1367); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1369 = 7'h3f == data1Frac_10 ? $signed(8'sh2e) : $signed(_GEN_1368); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1370 = 7'h40 == data1Frac_10 ? $signed(8'sh2d) : $signed(_GEN_1369); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1371 = 7'h41 == data1Frac_10 ? $signed(8'sh2d) : $signed(_GEN_1370); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1372 = 7'h42 == data1Frac_10 ? $signed(8'sh2d) : $signed(_GEN_1371); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1373 = 7'h43 == data1Frac_10 ? $signed(8'sh2d) : $signed(_GEN_1372); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1374 = 7'h44 == data1Frac_10 ? $signed(8'sh2c) : $signed(_GEN_1373); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1375 = 7'h45 == data1Frac_10 ? $signed(8'sh2c) : $signed(_GEN_1374); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1376 = 7'h46 == data1Frac_10 ? $signed(8'sh2c) : $signed(_GEN_1375); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1377 = 7'h47 == data1Frac_10 ? $signed(8'sh2c) : $signed(_GEN_1376); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1378 = 7'h48 == data1Frac_10 ? $signed(8'sh2b) : $signed(_GEN_1377); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1379 = 7'h49 == data1Frac_10 ? $signed(8'sh2b) : $signed(_GEN_1378); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1380 = 7'h4a == data1Frac_10 ? $signed(8'sh2b) : $signed(_GEN_1379); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1381 = 7'h4b == data1Frac_10 ? $signed(8'sh2b) : $signed(_GEN_1380); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1382 = 7'h4c == data1Frac_10 ? $signed(8'sh2a) : $signed(_GEN_1381); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1383 = 7'h4d == data1Frac_10 ? $signed(8'sh2a) : $signed(_GEN_1382); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1384 = 7'h4e == data1Frac_10 ? $signed(8'sh2a) : $signed(_GEN_1383); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1385 = 7'h4f == data1Frac_10 ? $signed(8'sh2a) : $signed(_GEN_1384); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1386 = 7'h50 == data1Frac_10 ? $signed(8'sh29) : $signed(_GEN_1385); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1387 = 7'h51 == data1Frac_10 ? $signed(8'sh29) : $signed(_GEN_1386); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1388 = 7'h52 == data1Frac_10 ? $signed(8'sh29) : $signed(_GEN_1387); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1389 = 7'h53 == data1Frac_10 ? $signed(8'sh29) : $signed(_GEN_1388); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1390 = 7'h54 == data1Frac_10 ? $signed(8'sh29) : $signed(_GEN_1389); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1391 = 7'h55 == data1Frac_10 ? $signed(8'sh28) : $signed(_GEN_1390); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1392 = 7'h56 == data1Frac_10 ? $signed(8'sh28) : $signed(_GEN_1391); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1393 = 7'h57 == data1Frac_10 ? $signed(8'sh28) : $signed(_GEN_1392); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1394 = 7'h58 == data1Frac_10 ? $signed(8'sh28) : $signed(_GEN_1393); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1395 = 7'h59 == data1Frac_10 ? $signed(8'sh28) : $signed(_GEN_1394); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1396 = 7'h5a == data1Frac_10 ? $signed(8'sh27) : $signed(_GEN_1395); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1397 = 7'h5b == data1Frac_10 ? $signed(8'sh27) : $signed(_GEN_1396); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1398 = 7'h5c == data1Frac_10 ? $signed(8'sh27) : $signed(_GEN_1397); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1399 = 7'h5d == data1Frac_10 ? $signed(8'sh27) : $signed(_GEN_1398); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1400 = 7'h5e == data1Frac_10 ? $signed(8'sh26) : $signed(_GEN_1399); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1401 = 7'h5f == data1Frac_10 ? $signed(8'sh26) : $signed(_GEN_1400); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1402 = 7'h60 == data1Frac_10 ? $signed(8'sh26) : $signed(_GEN_1401); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1403 = 7'h61 == data1Frac_10 ? $signed(8'sh26) : $signed(_GEN_1402); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1404 = 7'h62 == data1Frac_10 ? $signed(8'sh26) : $signed(_GEN_1403); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1405 = 7'h63 == data1Frac_10 ? $signed(8'sh25) : $signed(_GEN_1404); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1406 = 7'h64 == data1Frac_10 ? $signed(8'sh25) : $signed(_GEN_1405); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1407 = 7'h65 == data1Frac_10 ? $signed(8'sh25) : $signed(_GEN_1406); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1408 = 7'h66 == data1Frac_10 ? $signed(8'sh25) : $signed(_GEN_1407); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1409 = 7'h67 == data1Frac_10 ? $signed(8'sh25) : $signed(_GEN_1408); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1410 = 7'h68 == data1Frac_10 ? $signed(8'sh24) : $signed(_GEN_1409); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1411 = 7'h69 == data1Frac_10 ? $signed(8'sh24) : $signed(_GEN_1410); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1412 = 7'h6a == data1Frac_10 ? $signed(8'sh24) : $signed(_GEN_1411); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1413 = 7'h6b == data1Frac_10 ? $signed(8'sh24) : $signed(_GEN_1412); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1414 = 7'h6c == data1Frac_10 ? $signed(8'sh24) : $signed(_GEN_1413); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1415 = 7'h6d == data1Frac_10 ? $signed(8'sh23) : $signed(_GEN_1414); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1416 = 7'h6e == data1Frac_10 ? $signed(8'sh23) : $signed(_GEN_1415); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1417 = 7'h6f == data1Frac_10 ? $signed(8'sh23) : $signed(_GEN_1416); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1418 = 7'h70 == data1Frac_10 ? $signed(8'sh23) : $signed(_GEN_1417); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1419 = 7'h71 == data1Frac_10 ? $signed(8'sh23) : $signed(_GEN_1418); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1420 = 7'h72 == data1Frac_10 ? $signed(8'sh23) : $signed(_GEN_1419); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1421 = 7'h73 == data1Frac_10 ? $signed(8'sh22) : $signed(_GEN_1420); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1422 = 7'h74 == data1Frac_10 ? $signed(8'sh22) : $signed(_GEN_1421); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1423 = 7'h75 == data1Frac_10 ? $signed(8'sh22) : $signed(_GEN_1422); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1424 = 7'h76 == data1Frac_10 ? $signed(8'sh22) : $signed(_GEN_1423); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1425 = 7'h77 == data1Frac_10 ? $signed(8'sh22) : $signed(_GEN_1424); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1426 = 7'h78 == data1Frac_10 ? $signed(8'sh21) : $signed(_GEN_1425); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1427 = 7'h79 == data1Frac_10 ? $signed(8'sh21) : $signed(_GEN_1426); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1428 = 7'h7a == data1Frac_10 ? $signed(8'sh21) : $signed(_GEN_1427); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1429 = 7'h7b == data1Frac_10 ? $signed(8'sh21) : $signed(_GEN_1428); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1430 = 7'h7c == data1Frac_10 ? $signed(8'sh21) : $signed(_GEN_1429); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1431 = 7'h7d == data1Frac_10 ? $signed(8'sh21) : $signed(_GEN_1430); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1432 = 7'h7e == data1Frac_10 ? $signed(8'sh20) : $signed(_GEN_1431); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1433 = 7'h7f == data1Frac_10 ? $signed(8'sh20) : $signed(_GEN_1432); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_32 = $signed(_GEN_1433) >>> data1Int_10; // @[exponent.scala 38:85]
  reg [7:0] data2_10; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1437 = 7'h2 == data1Frac_11 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1438 = 7'h3 == data1Frac_11 ? $signed(8'sh3f) : $signed(_GEN_1437); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1439 = 7'h4 == data1Frac_11 ? $signed(8'sh3f) : $signed(_GEN_1438); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1440 = 7'h5 == data1Frac_11 ? $signed(8'sh3e) : $signed(_GEN_1439); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1441 = 7'h6 == data1Frac_11 ? $signed(8'sh3e) : $signed(_GEN_1440); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1442 = 7'h7 == data1Frac_11 ? $signed(8'sh3e) : $signed(_GEN_1441); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1443 = 7'h8 == data1Frac_11 ? $signed(8'sh3d) : $signed(_GEN_1442); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1444 = 7'h9 == data1Frac_11 ? $signed(8'sh3d) : $signed(_GEN_1443); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1445 = 7'ha == data1Frac_11 ? $signed(8'sh3d) : $signed(_GEN_1444); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1446 = 7'hb == data1Frac_11 ? $signed(8'sh3c) : $signed(_GEN_1445); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1447 = 7'hc == data1Frac_11 ? $signed(8'sh3c) : $signed(_GEN_1446); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1448 = 7'hd == data1Frac_11 ? $signed(8'sh3c) : $signed(_GEN_1447); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1449 = 7'he == data1Frac_11 ? $signed(8'sh3b) : $signed(_GEN_1448); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1450 = 7'hf == data1Frac_11 ? $signed(8'sh3b) : $signed(_GEN_1449); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1451 = 7'h10 == data1Frac_11 ? $signed(8'sh3b) : $signed(_GEN_1450); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1452 = 7'h11 == data1Frac_11 ? $signed(8'sh3a) : $signed(_GEN_1451); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1453 = 7'h12 == data1Frac_11 ? $signed(8'sh3a) : $signed(_GEN_1452); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1454 = 7'h13 == data1Frac_11 ? $signed(8'sh3a) : $signed(_GEN_1453); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1455 = 7'h14 == data1Frac_11 ? $signed(8'sh39) : $signed(_GEN_1454); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1456 = 7'h15 == data1Frac_11 ? $signed(8'sh39) : $signed(_GEN_1455); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1457 = 7'h16 == data1Frac_11 ? $signed(8'sh39) : $signed(_GEN_1456); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1458 = 7'h17 == data1Frac_11 ? $signed(8'sh39) : $signed(_GEN_1457); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1459 = 7'h18 == data1Frac_11 ? $signed(8'sh38) : $signed(_GEN_1458); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1460 = 7'h19 == data1Frac_11 ? $signed(8'sh38) : $signed(_GEN_1459); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1461 = 7'h1a == data1Frac_11 ? $signed(8'sh38) : $signed(_GEN_1460); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1462 = 7'h1b == data1Frac_11 ? $signed(8'sh37) : $signed(_GEN_1461); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1463 = 7'h1c == data1Frac_11 ? $signed(8'sh37) : $signed(_GEN_1462); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1464 = 7'h1d == data1Frac_11 ? $signed(8'sh37) : $signed(_GEN_1463); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1465 = 7'h1e == data1Frac_11 ? $signed(8'sh36) : $signed(_GEN_1464); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1466 = 7'h1f == data1Frac_11 ? $signed(8'sh36) : $signed(_GEN_1465); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1467 = 7'h20 == data1Frac_11 ? $signed(8'sh36) : $signed(_GEN_1466); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1468 = 7'h21 == data1Frac_11 ? $signed(8'sh36) : $signed(_GEN_1467); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1469 = 7'h22 == data1Frac_11 ? $signed(8'sh35) : $signed(_GEN_1468); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1470 = 7'h23 == data1Frac_11 ? $signed(8'sh35) : $signed(_GEN_1469); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1471 = 7'h24 == data1Frac_11 ? $signed(8'sh35) : $signed(_GEN_1470); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1472 = 7'h25 == data1Frac_11 ? $signed(8'sh34) : $signed(_GEN_1471); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1473 = 7'h26 == data1Frac_11 ? $signed(8'sh34) : $signed(_GEN_1472); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1474 = 7'h27 == data1Frac_11 ? $signed(8'sh34) : $signed(_GEN_1473); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1475 = 7'h28 == data1Frac_11 ? $signed(8'sh34) : $signed(_GEN_1474); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1476 = 7'h29 == data1Frac_11 ? $signed(8'sh33) : $signed(_GEN_1475); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1477 = 7'h2a == data1Frac_11 ? $signed(8'sh33) : $signed(_GEN_1476); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1478 = 7'h2b == data1Frac_11 ? $signed(8'sh33) : $signed(_GEN_1477); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1479 = 7'h2c == data1Frac_11 ? $signed(8'sh32) : $signed(_GEN_1478); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1480 = 7'h2d == data1Frac_11 ? $signed(8'sh32) : $signed(_GEN_1479); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1481 = 7'h2e == data1Frac_11 ? $signed(8'sh32) : $signed(_GEN_1480); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1482 = 7'h2f == data1Frac_11 ? $signed(8'sh32) : $signed(_GEN_1481); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1483 = 7'h30 == data1Frac_11 ? $signed(8'sh31) : $signed(_GEN_1482); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1484 = 7'h31 == data1Frac_11 ? $signed(8'sh31) : $signed(_GEN_1483); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1485 = 7'h32 == data1Frac_11 ? $signed(8'sh31) : $signed(_GEN_1484); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1486 = 7'h33 == data1Frac_11 ? $signed(8'sh31) : $signed(_GEN_1485); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1487 = 7'h34 == data1Frac_11 ? $signed(8'sh30) : $signed(_GEN_1486); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1488 = 7'h35 == data1Frac_11 ? $signed(8'sh30) : $signed(_GEN_1487); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1489 = 7'h36 == data1Frac_11 ? $signed(8'sh30) : $signed(_GEN_1488); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1490 = 7'h37 == data1Frac_11 ? $signed(8'sh30) : $signed(_GEN_1489); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1491 = 7'h38 == data1Frac_11 ? $signed(8'sh2f) : $signed(_GEN_1490); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1492 = 7'h39 == data1Frac_11 ? $signed(8'sh2f) : $signed(_GEN_1491); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1493 = 7'h3a == data1Frac_11 ? $signed(8'sh2f) : $signed(_GEN_1492); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1494 = 7'h3b == data1Frac_11 ? $signed(8'sh2e) : $signed(_GEN_1493); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1495 = 7'h3c == data1Frac_11 ? $signed(8'sh2e) : $signed(_GEN_1494); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1496 = 7'h3d == data1Frac_11 ? $signed(8'sh2e) : $signed(_GEN_1495); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1497 = 7'h3e == data1Frac_11 ? $signed(8'sh2e) : $signed(_GEN_1496); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1498 = 7'h3f == data1Frac_11 ? $signed(8'sh2e) : $signed(_GEN_1497); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1499 = 7'h40 == data1Frac_11 ? $signed(8'sh2d) : $signed(_GEN_1498); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1500 = 7'h41 == data1Frac_11 ? $signed(8'sh2d) : $signed(_GEN_1499); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1501 = 7'h42 == data1Frac_11 ? $signed(8'sh2d) : $signed(_GEN_1500); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1502 = 7'h43 == data1Frac_11 ? $signed(8'sh2d) : $signed(_GEN_1501); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1503 = 7'h44 == data1Frac_11 ? $signed(8'sh2c) : $signed(_GEN_1502); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1504 = 7'h45 == data1Frac_11 ? $signed(8'sh2c) : $signed(_GEN_1503); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1505 = 7'h46 == data1Frac_11 ? $signed(8'sh2c) : $signed(_GEN_1504); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1506 = 7'h47 == data1Frac_11 ? $signed(8'sh2c) : $signed(_GEN_1505); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1507 = 7'h48 == data1Frac_11 ? $signed(8'sh2b) : $signed(_GEN_1506); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1508 = 7'h49 == data1Frac_11 ? $signed(8'sh2b) : $signed(_GEN_1507); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1509 = 7'h4a == data1Frac_11 ? $signed(8'sh2b) : $signed(_GEN_1508); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1510 = 7'h4b == data1Frac_11 ? $signed(8'sh2b) : $signed(_GEN_1509); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1511 = 7'h4c == data1Frac_11 ? $signed(8'sh2a) : $signed(_GEN_1510); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1512 = 7'h4d == data1Frac_11 ? $signed(8'sh2a) : $signed(_GEN_1511); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1513 = 7'h4e == data1Frac_11 ? $signed(8'sh2a) : $signed(_GEN_1512); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1514 = 7'h4f == data1Frac_11 ? $signed(8'sh2a) : $signed(_GEN_1513); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1515 = 7'h50 == data1Frac_11 ? $signed(8'sh29) : $signed(_GEN_1514); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1516 = 7'h51 == data1Frac_11 ? $signed(8'sh29) : $signed(_GEN_1515); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1517 = 7'h52 == data1Frac_11 ? $signed(8'sh29) : $signed(_GEN_1516); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1518 = 7'h53 == data1Frac_11 ? $signed(8'sh29) : $signed(_GEN_1517); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1519 = 7'h54 == data1Frac_11 ? $signed(8'sh29) : $signed(_GEN_1518); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1520 = 7'h55 == data1Frac_11 ? $signed(8'sh28) : $signed(_GEN_1519); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1521 = 7'h56 == data1Frac_11 ? $signed(8'sh28) : $signed(_GEN_1520); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1522 = 7'h57 == data1Frac_11 ? $signed(8'sh28) : $signed(_GEN_1521); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1523 = 7'h58 == data1Frac_11 ? $signed(8'sh28) : $signed(_GEN_1522); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1524 = 7'h59 == data1Frac_11 ? $signed(8'sh28) : $signed(_GEN_1523); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1525 = 7'h5a == data1Frac_11 ? $signed(8'sh27) : $signed(_GEN_1524); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1526 = 7'h5b == data1Frac_11 ? $signed(8'sh27) : $signed(_GEN_1525); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1527 = 7'h5c == data1Frac_11 ? $signed(8'sh27) : $signed(_GEN_1526); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1528 = 7'h5d == data1Frac_11 ? $signed(8'sh27) : $signed(_GEN_1527); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1529 = 7'h5e == data1Frac_11 ? $signed(8'sh26) : $signed(_GEN_1528); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1530 = 7'h5f == data1Frac_11 ? $signed(8'sh26) : $signed(_GEN_1529); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1531 = 7'h60 == data1Frac_11 ? $signed(8'sh26) : $signed(_GEN_1530); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1532 = 7'h61 == data1Frac_11 ? $signed(8'sh26) : $signed(_GEN_1531); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1533 = 7'h62 == data1Frac_11 ? $signed(8'sh26) : $signed(_GEN_1532); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1534 = 7'h63 == data1Frac_11 ? $signed(8'sh25) : $signed(_GEN_1533); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1535 = 7'h64 == data1Frac_11 ? $signed(8'sh25) : $signed(_GEN_1534); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1536 = 7'h65 == data1Frac_11 ? $signed(8'sh25) : $signed(_GEN_1535); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1537 = 7'h66 == data1Frac_11 ? $signed(8'sh25) : $signed(_GEN_1536); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1538 = 7'h67 == data1Frac_11 ? $signed(8'sh25) : $signed(_GEN_1537); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1539 = 7'h68 == data1Frac_11 ? $signed(8'sh24) : $signed(_GEN_1538); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1540 = 7'h69 == data1Frac_11 ? $signed(8'sh24) : $signed(_GEN_1539); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1541 = 7'h6a == data1Frac_11 ? $signed(8'sh24) : $signed(_GEN_1540); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1542 = 7'h6b == data1Frac_11 ? $signed(8'sh24) : $signed(_GEN_1541); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1543 = 7'h6c == data1Frac_11 ? $signed(8'sh24) : $signed(_GEN_1542); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1544 = 7'h6d == data1Frac_11 ? $signed(8'sh23) : $signed(_GEN_1543); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1545 = 7'h6e == data1Frac_11 ? $signed(8'sh23) : $signed(_GEN_1544); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1546 = 7'h6f == data1Frac_11 ? $signed(8'sh23) : $signed(_GEN_1545); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1547 = 7'h70 == data1Frac_11 ? $signed(8'sh23) : $signed(_GEN_1546); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1548 = 7'h71 == data1Frac_11 ? $signed(8'sh23) : $signed(_GEN_1547); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1549 = 7'h72 == data1Frac_11 ? $signed(8'sh23) : $signed(_GEN_1548); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1550 = 7'h73 == data1Frac_11 ? $signed(8'sh22) : $signed(_GEN_1549); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1551 = 7'h74 == data1Frac_11 ? $signed(8'sh22) : $signed(_GEN_1550); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1552 = 7'h75 == data1Frac_11 ? $signed(8'sh22) : $signed(_GEN_1551); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1553 = 7'h76 == data1Frac_11 ? $signed(8'sh22) : $signed(_GEN_1552); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1554 = 7'h77 == data1Frac_11 ? $signed(8'sh22) : $signed(_GEN_1553); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1555 = 7'h78 == data1Frac_11 ? $signed(8'sh21) : $signed(_GEN_1554); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1556 = 7'h79 == data1Frac_11 ? $signed(8'sh21) : $signed(_GEN_1555); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1557 = 7'h7a == data1Frac_11 ? $signed(8'sh21) : $signed(_GEN_1556); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1558 = 7'h7b == data1Frac_11 ? $signed(8'sh21) : $signed(_GEN_1557); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1559 = 7'h7c == data1Frac_11 ? $signed(8'sh21) : $signed(_GEN_1558); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1560 = 7'h7d == data1Frac_11 ? $signed(8'sh21) : $signed(_GEN_1559); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1561 = 7'h7e == data1Frac_11 ? $signed(8'sh20) : $signed(_GEN_1560); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1562 = 7'h7f == data1Frac_11 ? $signed(8'sh20) : $signed(_GEN_1561); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_35 = $signed(_GEN_1562) >>> data1Int_11; // @[exponent.scala 38:85]
  reg [7:0] data2_11; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1566 = 7'h2 == data1Frac_12 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1567 = 7'h3 == data1Frac_12 ? $signed(8'sh3f) : $signed(_GEN_1566); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1568 = 7'h4 == data1Frac_12 ? $signed(8'sh3f) : $signed(_GEN_1567); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1569 = 7'h5 == data1Frac_12 ? $signed(8'sh3e) : $signed(_GEN_1568); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1570 = 7'h6 == data1Frac_12 ? $signed(8'sh3e) : $signed(_GEN_1569); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1571 = 7'h7 == data1Frac_12 ? $signed(8'sh3e) : $signed(_GEN_1570); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1572 = 7'h8 == data1Frac_12 ? $signed(8'sh3d) : $signed(_GEN_1571); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1573 = 7'h9 == data1Frac_12 ? $signed(8'sh3d) : $signed(_GEN_1572); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1574 = 7'ha == data1Frac_12 ? $signed(8'sh3d) : $signed(_GEN_1573); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1575 = 7'hb == data1Frac_12 ? $signed(8'sh3c) : $signed(_GEN_1574); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1576 = 7'hc == data1Frac_12 ? $signed(8'sh3c) : $signed(_GEN_1575); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1577 = 7'hd == data1Frac_12 ? $signed(8'sh3c) : $signed(_GEN_1576); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1578 = 7'he == data1Frac_12 ? $signed(8'sh3b) : $signed(_GEN_1577); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1579 = 7'hf == data1Frac_12 ? $signed(8'sh3b) : $signed(_GEN_1578); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1580 = 7'h10 == data1Frac_12 ? $signed(8'sh3b) : $signed(_GEN_1579); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1581 = 7'h11 == data1Frac_12 ? $signed(8'sh3a) : $signed(_GEN_1580); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1582 = 7'h12 == data1Frac_12 ? $signed(8'sh3a) : $signed(_GEN_1581); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1583 = 7'h13 == data1Frac_12 ? $signed(8'sh3a) : $signed(_GEN_1582); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1584 = 7'h14 == data1Frac_12 ? $signed(8'sh39) : $signed(_GEN_1583); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1585 = 7'h15 == data1Frac_12 ? $signed(8'sh39) : $signed(_GEN_1584); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1586 = 7'h16 == data1Frac_12 ? $signed(8'sh39) : $signed(_GEN_1585); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1587 = 7'h17 == data1Frac_12 ? $signed(8'sh39) : $signed(_GEN_1586); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1588 = 7'h18 == data1Frac_12 ? $signed(8'sh38) : $signed(_GEN_1587); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1589 = 7'h19 == data1Frac_12 ? $signed(8'sh38) : $signed(_GEN_1588); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1590 = 7'h1a == data1Frac_12 ? $signed(8'sh38) : $signed(_GEN_1589); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1591 = 7'h1b == data1Frac_12 ? $signed(8'sh37) : $signed(_GEN_1590); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1592 = 7'h1c == data1Frac_12 ? $signed(8'sh37) : $signed(_GEN_1591); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1593 = 7'h1d == data1Frac_12 ? $signed(8'sh37) : $signed(_GEN_1592); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1594 = 7'h1e == data1Frac_12 ? $signed(8'sh36) : $signed(_GEN_1593); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1595 = 7'h1f == data1Frac_12 ? $signed(8'sh36) : $signed(_GEN_1594); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1596 = 7'h20 == data1Frac_12 ? $signed(8'sh36) : $signed(_GEN_1595); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1597 = 7'h21 == data1Frac_12 ? $signed(8'sh36) : $signed(_GEN_1596); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1598 = 7'h22 == data1Frac_12 ? $signed(8'sh35) : $signed(_GEN_1597); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1599 = 7'h23 == data1Frac_12 ? $signed(8'sh35) : $signed(_GEN_1598); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1600 = 7'h24 == data1Frac_12 ? $signed(8'sh35) : $signed(_GEN_1599); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1601 = 7'h25 == data1Frac_12 ? $signed(8'sh34) : $signed(_GEN_1600); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1602 = 7'h26 == data1Frac_12 ? $signed(8'sh34) : $signed(_GEN_1601); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1603 = 7'h27 == data1Frac_12 ? $signed(8'sh34) : $signed(_GEN_1602); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1604 = 7'h28 == data1Frac_12 ? $signed(8'sh34) : $signed(_GEN_1603); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1605 = 7'h29 == data1Frac_12 ? $signed(8'sh33) : $signed(_GEN_1604); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1606 = 7'h2a == data1Frac_12 ? $signed(8'sh33) : $signed(_GEN_1605); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1607 = 7'h2b == data1Frac_12 ? $signed(8'sh33) : $signed(_GEN_1606); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1608 = 7'h2c == data1Frac_12 ? $signed(8'sh32) : $signed(_GEN_1607); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1609 = 7'h2d == data1Frac_12 ? $signed(8'sh32) : $signed(_GEN_1608); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1610 = 7'h2e == data1Frac_12 ? $signed(8'sh32) : $signed(_GEN_1609); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1611 = 7'h2f == data1Frac_12 ? $signed(8'sh32) : $signed(_GEN_1610); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1612 = 7'h30 == data1Frac_12 ? $signed(8'sh31) : $signed(_GEN_1611); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1613 = 7'h31 == data1Frac_12 ? $signed(8'sh31) : $signed(_GEN_1612); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1614 = 7'h32 == data1Frac_12 ? $signed(8'sh31) : $signed(_GEN_1613); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1615 = 7'h33 == data1Frac_12 ? $signed(8'sh31) : $signed(_GEN_1614); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1616 = 7'h34 == data1Frac_12 ? $signed(8'sh30) : $signed(_GEN_1615); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1617 = 7'h35 == data1Frac_12 ? $signed(8'sh30) : $signed(_GEN_1616); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1618 = 7'h36 == data1Frac_12 ? $signed(8'sh30) : $signed(_GEN_1617); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1619 = 7'h37 == data1Frac_12 ? $signed(8'sh30) : $signed(_GEN_1618); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1620 = 7'h38 == data1Frac_12 ? $signed(8'sh2f) : $signed(_GEN_1619); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1621 = 7'h39 == data1Frac_12 ? $signed(8'sh2f) : $signed(_GEN_1620); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1622 = 7'h3a == data1Frac_12 ? $signed(8'sh2f) : $signed(_GEN_1621); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1623 = 7'h3b == data1Frac_12 ? $signed(8'sh2e) : $signed(_GEN_1622); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1624 = 7'h3c == data1Frac_12 ? $signed(8'sh2e) : $signed(_GEN_1623); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1625 = 7'h3d == data1Frac_12 ? $signed(8'sh2e) : $signed(_GEN_1624); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1626 = 7'h3e == data1Frac_12 ? $signed(8'sh2e) : $signed(_GEN_1625); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1627 = 7'h3f == data1Frac_12 ? $signed(8'sh2e) : $signed(_GEN_1626); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1628 = 7'h40 == data1Frac_12 ? $signed(8'sh2d) : $signed(_GEN_1627); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1629 = 7'h41 == data1Frac_12 ? $signed(8'sh2d) : $signed(_GEN_1628); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1630 = 7'h42 == data1Frac_12 ? $signed(8'sh2d) : $signed(_GEN_1629); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1631 = 7'h43 == data1Frac_12 ? $signed(8'sh2d) : $signed(_GEN_1630); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1632 = 7'h44 == data1Frac_12 ? $signed(8'sh2c) : $signed(_GEN_1631); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1633 = 7'h45 == data1Frac_12 ? $signed(8'sh2c) : $signed(_GEN_1632); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1634 = 7'h46 == data1Frac_12 ? $signed(8'sh2c) : $signed(_GEN_1633); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1635 = 7'h47 == data1Frac_12 ? $signed(8'sh2c) : $signed(_GEN_1634); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1636 = 7'h48 == data1Frac_12 ? $signed(8'sh2b) : $signed(_GEN_1635); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1637 = 7'h49 == data1Frac_12 ? $signed(8'sh2b) : $signed(_GEN_1636); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1638 = 7'h4a == data1Frac_12 ? $signed(8'sh2b) : $signed(_GEN_1637); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1639 = 7'h4b == data1Frac_12 ? $signed(8'sh2b) : $signed(_GEN_1638); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1640 = 7'h4c == data1Frac_12 ? $signed(8'sh2a) : $signed(_GEN_1639); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1641 = 7'h4d == data1Frac_12 ? $signed(8'sh2a) : $signed(_GEN_1640); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1642 = 7'h4e == data1Frac_12 ? $signed(8'sh2a) : $signed(_GEN_1641); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1643 = 7'h4f == data1Frac_12 ? $signed(8'sh2a) : $signed(_GEN_1642); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1644 = 7'h50 == data1Frac_12 ? $signed(8'sh29) : $signed(_GEN_1643); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1645 = 7'h51 == data1Frac_12 ? $signed(8'sh29) : $signed(_GEN_1644); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1646 = 7'h52 == data1Frac_12 ? $signed(8'sh29) : $signed(_GEN_1645); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1647 = 7'h53 == data1Frac_12 ? $signed(8'sh29) : $signed(_GEN_1646); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1648 = 7'h54 == data1Frac_12 ? $signed(8'sh29) : $signed(_GEN_1647); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1649 = 7'h55 == data1Frac_12 ? $signed(8'sh28) : $signed(_GEN_1648); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1650 = 7'h56 == data1Frac_12 ? $signed(8'sh28) : $signed(_GEN_1649); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1651 = 7'h57 == data1Frac_12 ? $signed(8'sh28) : $signed(_GEN_1650); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1652 = 7'h58 == data1Frac_12 ? $signed(8'sh28) : $signed(_GEN_1651); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1653 = 7'h59 == data1Frac_12 ? $signed(8'sh28) : $signed(_GEN_1652); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1654 = 7'h5a == data1Frac_12 ? $signed(8'sh27) : $signed(_GEN_1653); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1655 = 7'h5b == data1Frac_12 ? $signed(8'sh27) : $signed(_GEN_1654); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1656 = 7'h5c == data1Frac_12 ? $signed(8'sh27) : $signed(_GEN_1655); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1657 = 7'h5d == data1Frac_12 ? $signed(8'sh27) : $signed(_GEN_1656); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1658 = 7'h5e == data1Frac_12 ? $signed(8'sh26) : $signed(_GEN_1657); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1659 = 7'h5f == data1Frac_12 ? $signed(8'sh26) : $signed(_GEN_1658); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1660 = 7'h60 == data1Frac_12 ? $signed(8'sh26) : $signed(_GEN_1659); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1661 = 7'h61 == data1Frac_12 ? $signed(8'sh26) : $signed(_GEN_1660); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1662 = 7'h62 == data1Frac_12 ? $signed(8'sh26) : $signed(_GEN_1661); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1663 = 7'h63 == data1Frac_12 ? $signed(8'sh25) : $signed(_GEN_1662); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1664 = 7'h64 == data1Frac_12 ? $signed(8'sh25) : $signed(_GEN_1663); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1665 = 7'h65 == data1Frac_12 ? $signed(8'sh25) : $signed(_GEN_1664); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1666 = 7'h66 == data1Frac_12 ? $signed(8'sh25) : $signed(_GEN_1665); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1667 = 7'h67 == data1Frac_12 ? $signed(8'sh25) : $signed(_GEN_1666); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1668 = 7'h68 == data1Frac_12 ? $signed(8'sh24) : $signed(_GEN_1667); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1669 = 7'h69 == data1Frac_12 ? $signed(8'sh24) : $signed(_GEN_1668); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1670 = 7'h6a == data1Frac_12 ? $signed(8'sh24) : $signed(_GEN_1669); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1671 = 7'h6b == data1Frac_12 ? $signed(8'sh24) : $signed(_GEN_1670); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1672 = 7'h6c == data1Frac_12 ? $signed(8'sh24) : $signed(_GEN_1671); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1673 = 7'h6d == data1Frac_12 ? $signed(8'sh23) : $signed(_GEN_1672); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1674 = 7'h6e == data1Frac_12 ? $signed(8'sh23) : $signed(_GEN_1673); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1675 = 7'h6f == data1Frac_12 ? $signed(8'sh23) : $signed(_GEN_1674); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1676 = 7'h70 == data1Frac_12 ? $signed(8'sh23) : $signed(_GEN_1675); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1677 = 7'h71 == data1Frac_12 ? $signed(8'sh23) : $signed(_GEN_1676); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1678 = 7'h72 == data1Frac_12 ? $signed(8'sh23) : $signed(_GEN_1677); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1679 = 7'h73 == data1Frac_12 ? $signed(8'sh22) : $signed(_GEN_1678); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1680 = 7'h74 == data1Frac_12 ? $signed(8'sh22) : $signed(_GEN_1679); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1681 = 7'h75 == data1Frac_12 ? $signed(8'sh22) : $signed(_GEN_1680); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1682 = 7'h76 == data1Frac_12 ? $signed(8'sh22) : $signed(_GEN_1681); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1683 = 7'h77 == data1Frac_12 ? $signed(8'sh22) : $signed(_GEN_1682); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1684 = 7'h78 == data1Frac_12 ? $signed(8'sh21) : $signed(_GEN_1683); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1685 = 7'h79 == data1Frac_12 ? $signed(8'sh21) : $signed(_GEN_1684); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1686 = 7'h7a == data1Frac_12 ? $signed(8'sh21) : $signed(_GEN_1685); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1687 = 7'h7b == data1Frac_12 ? $signed(8'sh21) : $signed(_GEN_1686); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1688 = 7'h7c == data1Frac_12 ? $signed(8'sh21) : $signed(_GEN_1687); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1689 = 7'h7d == data1Frac_12 ? $signed(8'sh21) : $signed(_GEN_1688); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1690 = 7'h7e == data1Frac_12 ? $signed(8'sh20) : $signed(_GEN_1689); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1691 = 7'h7f == data1Frac_12 ? $signed(8'sh20) : $signed(_GEN_1690); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_38 = $signed(_GEN_1691) >>> data1Int_12; // @[exponent.scala 38:85]
  reg [7:0] data2_12; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1695 = 7'h2 == data1Frac_13 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1696 = 7'h3 == data1Frac_13 ? $signed(8'sh3f) : $signed(_GEN_1695); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1697 = 7'h4 == data1Frac_13 ? $signed(8'sh3f) : $signed(_GEN_1696); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1698 = 7'h5 == data1Frac_13 ? $signed(8'sh3e) : $signed(_GEN_1697); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1699 = 7'h6 == data1Frac_13 ? $signed(8'sh3e) : $signed(_GEN_1698); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1700 = 7'h7 == data1Frac_13 ? $signed(8'sh3e) : $signed(_GEN_1699); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1701 = 7'h8 == data1Frac_13 ? $signed(8'sh3d) : $signed(_GEN_1700); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1702 = 7'h9 == data1Frac_13 ? $signed(8'sh3d) : $signed(_GEN_1701); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1703 = 7'ha == data1Frac_13 ? $signed(8'sh3d) : $signed(_GEN_1702); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1704 = 7'hb == data1Frac_13 ? $signed(8'sh3c) : $signed(_GEN_1703); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1705 = 7'hc == data1Frac_13 ? $signed(8'sh3c) : $signed(_GEN_1704); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1706 = 7'hd == data1Frac_13 ? $signed(8'sh3c) : $signed(_GEN_1705); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1707 = 7'he == data1Frac_13 ? $signed(8'sh3b) : $signed(_GEN_1706); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1708 = 7'hf == data1Frac_13 ? $signed(8'sh3b) : $signed(_GEN_1707); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1709 = 7'h10 == data1Frac_13 ? $signed(8'sh3b) : $signed(_GEN_1708); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1710 = 7'h11 == data1Frac_13 ? $signed(8'sh3a) : $signed(_GEN_1709); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1711 = 7'h12 == data1Frac_13 ? $signed(8'sh3a) : $signed(_GEN_1710); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1712 = 7'h13 == data1Frac_13 ? $signed(8'sh3a) : $signed(_GEN_1711); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1713 = 7'h14 == data1Frac_13 ? $signed(8'sh39) : $signed(_GEN_1712); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1714 = 7'h15 == data1Frac_13 ? $signed(8'sh39) : $signed(_GEN_1713); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1715 = 7'h16 == data1Frac_13 ? $signed(8'sh39) : $signed(_GEN_1714); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1716 = 7'h17 == data1Frac_13 ? $signed(8'sh39) : $signed(_GEN_1715); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1717 = 7'h18 == data1Frac_13 ? $signed(8'sh38) : $signed(_GEN_1716); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1718 = 7'h19 == data1Frac_13 ? $signed(8'sh38) : $signed(_GEN_1717); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1719 = 7'h1a == data1Frac_13 ? $signed(8'sh38) : $signed(_GEN_1718); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1720 = 7'h1b == data1Frac_13 ? $signed(8'sh37) : $signed(_GEN_1719); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1721 = 7'h1c == data1Frac_13 ? $signed(8'sh37) : $signed(_GEN_1720); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1722 = 7'h1d == data1Frac_13 ? $signed(8'sh37) : $signed(_GEN_1721); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1723 = 7'h1e == data1Frac_13 ? $signed(8'sh36) : $signed(_GEN_1722); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1724 = 7'h1f == data1Frac_13 ? $signed(8'sh36) : $signed(_GEN_1723); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1725 = 7'h20 == data1Frac_13 ? $signed(8'sh36) : $signed(_GEN_1724); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1726 = 7'h21 == data1Frac_13 ? $signed(8'sh36) : $signed(_GEN_1725); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1727 = 7'h22 == data1Frac_13 ? $signed(8'sh35) : $signed(_GEN_1726); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1728 = 7'h23 == data1Frac_13 ? $signed(8'sh35) : $signed(_GEN_1727); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1729 = 7'h24 == data1Frac_13 ? $signed(8'sh35) : $signed(_GEN_1728); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1730 = 7'h25 == data1Frac_13 ? $signed(8'sh34) : $signed(_GEN_1729); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1731 = 7'h26 == data1Frac_13 ? $signed(8'sh34) : $signed(_GEN_1730); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1732 = 7'h27 == data1Frac_13 ? $signed(8'sh34) : $signed(_GEN_1731); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1733 = 7'h28 == data1Frac_13 ? $signed(8'sh34) : $signed(_GEN_1732); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1734 = 7'h29 == data1Frac_13 ? $signed(8'sh33) : $signed(_GEN_1733); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1735 = 7'h2a == data1Frac_13 ? $signed(8'sh33) : $signed(_GEN_1734); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1736 = 7'h2b == data1Frac_13 ? $signed(8'sh33) : $signed(_GEN_1735); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1737 = 7'h2c == data1Frac_13 ? $signed(8'sh32) : $signed(_GEN_1736); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1738 = 7'h2d == data1Frac_13 ? $signed(8'sh32) : $signed(_GEN_1737); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1739 = 7'h2e == data1Frac_13 ? $signed(8'sh32) : $signed(_GEN_1738); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1740 = 7'h2f == data1Frac_13 ? $signed(8'sh32) : $signed(_GEN_1739); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1741 = 7'h30 == data1Frac_13 ? $signed(8'sh31) : $signed(_GEN_1740); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1742 = 7'h31 == data1Frac_13 ? $signed(8'sh31) : $signed(_GEN_1741); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1743 = 7'h32 == data1Frac_13 ? $signed(8'sh31) : $signed(_GEN_1742); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1744 = 7'h33 == data1Frac_13 ? $signed(8'sh31) : $signed(_GEN_1743); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1745 = 7'h34 == data1Frac_13 ? $signed(8'sh30) : $signed(_GEN_1744); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1746 = 7'h35 == data1Frac_13 ? $signed(8'sh30) : $signed(_GEN_1745); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1747 = 7'h36 == data1Frac_13 ? $signed(8'sh30) : $signed(_GEN_1746); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1748 = 7'h37 == data1Frac_13 ? $signed(8'sh30) : $signed(_GEN_1747); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1749 = 7'h38 == data1Frac_13 ? $signed(8'sh2f) : $signed(_GEN_1748); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1750 = 7'h39 == data1Frac_13 ? $signed(8'sh2f) : $signed(_GEN_1749); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1751 = 7'h3a == data1Frac_13 ? $signed(8'sh2f) : $signed(_GEN_1750); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1752 = 7'h3b == data1Frac_13 ? $signed(8'sh2e) : $signed(_GEN_1751); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1753 = 7'h3c == data1Frac_13 ? $signed(8'sh2e) : $signed(_GEN_1752); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1754 = 7'h3d == data1Frac_13 ? $signed(8'sh2e) : $signed(_GEN_1753); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1755 = 7'h3e == data1Frac_13 ? $signed(8'sh2e) : $signed(_GEN_1754); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1756 = 7'h3f == data1Frac_13 ? $signed(8'sh2e) : $signed(_GEN_1755); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1757 = 7'h40 == data1Frac_13 ? $signed(8'sh2d) : $signed(_GEN_1756); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1758 = 7'h41 == data1Frac_13 ? $signed(8'sh2d) : $signed(_GEN_1757); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1759 = 7'h42 == data1Frac_13 ? $signed(8'sh2d) : $signed(_GEN_1758); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1760 = 7'h43 == data1Frac_13 ? $signed(8'sh2d) : $signed(_GEN_1759); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1761 = 7'h44 == data1Frac_13 ? $signed(8'sh2c) : $signed(_GEN_1760); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1762 = 7'h45 == data1Frac_13 ? $signed(8'sh2c) : $signed(_GEN_1761); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1763 = 7'h46 == data1Frac_13 ? $signed(8'sh2c) : $signed(_GEN_1762); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1764 = 7'h47 == data1Frac_13 ? $signed(8'sh2c) : $signed(_GEN_1763); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1765 = 7'h48 == data1Frac_13 ? $signed(8'sh2b) : $signed(_GEN_1764); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1766 = 7'h49 == data1Frac_13 ? $signed(8'sh2b) : $signed(_GEN_1765); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1767 = 7'h4a == data1Frac_13 ? $signed(8'sh2b) : $signed(_GEN_1766); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1768 = 7'h4b == data1Frac_13 ? $signed(8'sh2b) : $signed(_GEN_1767); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1769 = 7'h4c == data1Frac_13 ? $signed(8'sh2a) : $signed(_GEN_1768); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1770 = 7'h4d == data1Frac_13 ? $signed(8'sh2a) : $signed(_GEN_1769); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1771 = 7'h4e == data1Frac_13 ? $signed(8'sh2a) : $signed(_GEN_1770); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1772 = 7'h4f == data1Frac_13 ? $signed(8'sh2a) : $signed(_GEN_1771); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1773 = 7'h50 == data1Frac_13 ? $signed(8'sh29) : $signed(_GEN_1772); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1774 = 7'h51 == data1Frac_13 ? $signed(8'sh29) : $signed(_GEN_1773); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1775 = 7'h52 == data1Frac_13 ? $signed(8'sh29) : $signed(_GEN_1774); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1776 = 7'h53 == data1Frac_13 ? $signed(8'sh29) : $signed(_GEN_1775); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1777 = 7'h54 == data1Frac_13 ? $signed(8'sh29) : $signed(_GEN_1776); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1778 = 7'h55 == data1Frac_13 ? $signed(8'sh28) : $signed(_GEN_1777); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1779 = 7'h56 == data1Frac_13 ? $signed(8'sh28) : $signed(_GEN_1778); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1780 = 7'h57 == data1Frac_13 ? $signed(8'sh28) : $signed(_GEN_1779); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1781 = 7'h58 == data1Frac_13 ? $signed(8'sh28) : $signed(_GEN_1780); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1782 = 7'h59 == data1Frac_13 ? $signed(8'sh28) : $signed(_GEN_1781); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1783 = 7'h5a == data1Frac_13 ? $signed(8'sh27) : $signed(_GEN_1782); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1784 = 7'h5b == data1Frac_13 ? $signed(8'sh27) : $signed(_GEN_1783); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1785 = 7'h5c == data1Frac_13 ? $signed(8'sh27) : $signed(_GEN_1784); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1786 = 7'h5d == data1Frac_13 ? $signed(8'sh27) : $signed(_GEN_1785); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1787 = 7'h5e == data1Frac_13 ? $signed(8'sh26) : $signed(_GEN_1786); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1788 = 7'h5f == data1Frac_13 ? $signed(8'sh26) : $signed(_GEN_1787); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1789 = 7'h60 == data1Frac_13 ? $signed(8'sh26) : $signed(_GEN_1788); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1790 = 7'h61 == data1Frac_13 ? $signed(8'sh26) : $signed(_GEN_1789); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1791 = 7'h62 == data1Frac_13 ? $signed(8'sh26) : $signed(_GEN_1790); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1792 = 7'h63 == data1Frac_13 ? $signed(8'sh25) : $signed(_GEN_1791); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1793 = 7'h64 == data1Frac_13 ? $signed(8'sh25) : $signed(_GEN_1792); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1794 = 7'h65 == data1Frac_13 ? $signed(8'sh25) : $signed(_GEN_1793); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1795 = 7'h66 == data1Frac_13 ? $signed(8'sh25) : $signed(_GEN_1794); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1796 = 7'h67 == data1Frac_13 ? $signed(8'sh25) : $signed(_GEN_1795); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1797 = 7'h68 == data1Frac_13 ? $signed(8'sh24) : $signed(_GEN_1796); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1798 = 7'h69 == data1Frac_13 ? $signed(8'sh24) : $signed(_GEN_1797); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1799 = 7'h6a == data1Frac_13 ? $signed(8'sh24) : $signed(_GEN_1798); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1800 = 7'h6b == data1Frac_13 ? $signed(8'sh24) : $signed(_GEN_1799); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1801 = 7'h6c == data1Frac_13 ? $signed(8'sh24) : $signed(_GEN_1800); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1802 = 7'h6d == data1Frac_13 ? $signed(8'sh23) : $signed(_GEN_1801); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1803 = 7'h6e == data1Frac_13 ? $signed(8'sh23) : $signed(_GEN_1802); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1804 = 7'h6f == data1Frac_13 ? $signed(8'sh23) : $signed(_GEN_1803); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1805 = 7'h70 == data1Frac_13 ? $signed(8'sh23) : $signed(_GEN_1804); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1806 = 7'h71 == data1Frac_13 ? $signed(8'sh23) : $signed(_GEN_1805); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1807 = 7'h72 == data1Frac_13 ? $signed(8'sh23) : $signed(_GEN_1806); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1808 = 7'h73 == data1Frac_13 ? $signed(8'sh22) : $signed(_GEN_1807); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1809 = 7'h74 == data1Frac_13 ? $signed(8'sh22) : $signed(_GEN_1808); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1810 = 7'h75 == data1Frac_13 ? $signed(8'sh22) : $signed(_GEN_1809); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1811 = 7'h76 == data1Frac_13 ? $signed(8'sh22) : $signed(_GEN_1810); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1812 = 7'h77 == data1Frac_13 ? $signed(8'sh22) : $signed(_GEN_1811); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1813 = 7'h78 == data1Frac_13 ? $signed(8'sh21) : $signed(_GEN_1812); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1814 = 7'h79 == data1Frac_13 ? $signed(8'sh21) : $signed(_GEN_1813); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1815 = 7'h7a == data1Frac_13 ? $signed(8'sh21) : $signed(_GEN_1814); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1816 = 7'h7b == data1Frac_13 ? $signed(8'sh21) : $signed(_GEN_1815); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1817 = 7'h7c == data1Frac_13 ? $signed(8'sh21) : $signed(_GEN_1816); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1818 = 7'h7d == data1Frac_13 ? $signed(8'sh21) : $signed(_GEN_1817); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1819 = 7'h7e == data1Frac_13 ? $signed(8'sh20) : $signed(_GEN_1818); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1820 = 7'h7f == data1Frac_13 ? $signed(8'sh20) : $signed(_GEN_1819); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_41 = $signed(_GEN_1820) >>> data1Int_13; // @[exponent.scala 38:85]
  reg [7:0] data2_13; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1824 = 7'h2 == data1Frac_14 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1825 = 7'h3 == data1Frac_14 ? $signed(8'sh3f) : $signed(_GEN_1824); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1826 = 7'h4 == data1Frac_14 ? $signed(8'sh3f) : $signed(_GEN_1825); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1827 = 7'h5 == data1Frac_14 ? $signed(8'sh3e) : $signed(_GEN_1826); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1828 = 7'h6 == data1Frac_14 ? $signed(8'sh3e) : $signed(_GEN_1827); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1829 = 7'h7 == data1Frac_14 ? $signed(8'sh3e) : $signed(_GEN_1828); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1830 = 7'h8 == data1Frac_14 ? $signed(8'sh3d) : $signed(_GEN_1829); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1831 = 7'h9 == data1Frac_14 ? $signed(8'sh3d) : $signed(_GEN_1830); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1832 = 7'ha == data1Frac_14 ? $signed(8'sh3d) : $signed(_GEN_1831); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1833 = 7'hb == data1Frac_14 ? $signed(8'sh3c) : $signed(_GEN_1832); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1834 = 7'hc == data1Frac_14 ? $signed(8'sh3c) : $signed(_GEN_1833); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1835 = 7'hd == data1Frac_14 ? $signed(8'sh3c) : $signed(_GEN_1834); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1836 = 7'he == data1Frac_14 ? $signed(8'sh3b) : $signed(_GEN_1835); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1837 = 7'hf == data1Frac_14 ? $signed(8'sh3b) : $signed(_GEN_1836); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1838 = 7'h10 == data1Frac_14 ? $signed(8'sh3b) : $signed(_GEN_1837); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1839 = 7'h11 == data1Frac_14 ? $signed(8'sh3a) : $signed(_GEN_1838); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1840 = 7'h12 == data1Frac_14 ? $signed(8'sh3a) : $signed(_GEN_1839); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1841 = 7'h13 == data1Frac_14 ? $signed(8'sh3a) : $signed(_GEN_1840); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1842 = 7'h14 == data1Frac_14 ? $signed(8'sh39) : $signed(_GEN_1841); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1843 = 7'h15 == data1Frac_14 ? $signed(8'sh39) : $signed(_GEN_1842); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1844 = 7'h16 == data1Frac_14 ? $signed(8'sh39) : $signed(_GEN_1843); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1845 = 7'h17 == data1Frac_14 ? $signed(8'sh39) : $signed(_GEN_1844); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1846 = 7'h18 == data1Frac_14 ? $signed(8'sh38) : $signed(_GEN_1845); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1847 = 7'h19 == data1Frac_14 ? $signed(8'sh38) : $signed(_GEN_1846); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1848 = 7'h1a == data1Frac_14 ? $signed(8'sh38) : $signed(_GEN_1847); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1849 = 7'h1b == data1Frac_14 ? $signed(8'sh37) : $signed(_GEN_1848); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1850 = 7'h1c == data1Frac_14 ? $signed(8'sh37) : $signed(_GEN_1849); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1851 = 7'h1d == data1Frac_14 ? $signed(8'sh37) : $signed(_GEN_1850); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1852 = 7'h1e == data1Frac_14 ? $signed(8'sh36) : $signed(_GEN_1851); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1853 = 7'h1f == data1Frac_14 ? $signed(8'sh36) : $signed(_GEN_1852); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1854 = 7'h20 == data1Frac_14 ? $signed(8'sh36) : $signed(_GEN_1853); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1855 = 7'h21 == data1Frac_14 ? $signed(8'sh36) : $signed(_GEN_1854); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1856 = 7'h22 == data1Frac_14 ? $signed(8'sh35) : $signed(_GEN_1855); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1857 = 7'h23 == data1Frac_14 ? $signed(8'sh35) : $signed(_GEN_1856); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1858 = 7'h24 == data1Frac_14 ? $signed(8'sh35) : $signed(_GEN_1857); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1859 = 7'h25 == data1Frac_14 ? $signed(8'sh34) : $signed(_GEN_1858); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1860 = 7'h26 == data1Frac_14 ? $signed(8'sh34) : $signed(_GEN_1859); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1861 = 7'h27 == data1Frac_14 ? $signed(8'sh34) : $signed(_GEN_1860); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1862 = 7'h28 == data1Frac_14 ? $signed(8'sh34) : $signed(_GEN_1861); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1863 = 7'h29 == data1Frac_14 ? $signed(8'sh33) : $signed(_GEN_1862); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1864 = 7'h2a == data1Frac_14 ? $signed(8'sh33) : $signed(_GEN_1863); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1865 = 7'h2b == data1Frac_14 ? $signed(8'sh33) : $signed(_GEN_1864); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1866 = 7'h2c == data1Frac_14 ? $signed(8'sh32) : $signed(_GEN_1865); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1867 = 7'h2d == data1Frac_14 ? $signed(8'sh32) : $signed(_GEN_1866); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1868 = 7'h2e == data1Frac_14 ? $signed(8'sh32) : $signed(_GEN_1867); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1869 = 7'h2f == data1Frac_14 ? $signed(8'sh32) : $signed(_GEN_1868); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1870 = 7'h30 == data1Frac_14 ? $signed(8'sh31) : $signed(_GEN_1869); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1871 = 7'h31 == data1Frac_14 ? $signed(8'sh31) : $signed(_GEN_1870); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1872 = 7'h32 == data1Frac_14 ? $signed(8'sh31) : $signed(_GEN_1871); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1873 = 7'h33 == data1Frac_14 ? $signed(8'sh31) : $signed(_GEN_1872); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1874 = 7'h34 == data1Frac_14 ? $signed(8'sh30) : $signed(_GEN_1873); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1875 = 7'h35 == data1Frac_14 ? $signed(8'sh30) : $signed(_GEN_1874); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1876 = 7'h36 == data1Frac_14 ? $signed(8'sh30) : $signed(_GEN_1875); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1877 = 7'h37 == data1Frac_14 ? $signed(8'sh30) : $signed(_GEN_1876); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1878 = 7'h38 == data1Frac_14 ? $signed(8'sh2f) : $signed(_GEN_1877); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1879 = 7'h39 == data1Frac_14 ? $signed(8'sh2f) : $signed(_GEN_1878); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1880 = 7'h3a == data1Frac_14 ? $signed(8'sh2f) : $signed(_GEN_1879); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1881 = 7'h3b == data1Frac_14 ? $signed(8'sh2e) : $signed(_GEN_1880); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1882 = 7'h3c == data1Frac_14 ? $signed(8'sh2e) : $signed(_GEN_1881); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1883 = 7'h3d == data1Frac_14 ? $signed(8'sh2e) : $signed(_GEN_1882); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1884 = 7'h3e == data1Frac_14 ? $signed(8'sh2e) : $signed(_GEN_1883); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1885 = 7'h3f == data1Frac_14 ? $signed(8'sh2e) : $signed(_GEN_1884); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1886 = 7'h40 == data1Frac_14 ? $signed(8'sh2d) : $signed(_GEN_1885); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1887 = 7'h41 == data1Frac_14 ? $signed(8'sh2d) : $signed(_GEN_1886); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1888 = 7'h42 == data1Frac_14 ? $signed(8'sh2d) : $signed(_GEN_1887); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1889 = 7'h43 == data1Frac_14 ? $signed(8'sh2d) : $signed(_GEN_1888); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1890 = 7'h44 == data1Frac_14 ? $signed(8'sh2c) : $signed(_GEN_1889); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1891 = 7'h45 == data1Frac_14 ? $signed(8'sh2c) : $signed(_GEN_1890); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1892 = 7'h46 == data1Frac_14 ? $signed(8'sh2c) : $signed(_GEN_1891); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1893 = 7'h47 == data1Frac_14 ? $signed(8'sh2c) : $signed(_GEN_1892); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1894 = 7'h48 == data1Frac_14 ? $signed(8'sh2b) : $signed(_GEN_1893); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1895 = 7'h49 == data1Frac_14 ? $signed(8'sh2b) : $signed(_GEN_1894); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1896 = 7'h4a == data1Frac_14 ? $signed(8'sh2b) : $signed(_GEN_1895); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1897 = 7'h4b == data1Frac_14 ? $signed(8'sh2b) : $signed(_GEN_1896); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1898 = 7'h4c == data1Frac_14 ? $signed(8'sh2a) : $signed(_GEN_1897); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1899 = 7'h4d == data1Frac_14 ? $signed(8'sh2a) : $signed(_GEN_1898); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1900 = 7'h4e == data1Frac_14 ? $signed(8'sh2a) : $signed(_GEN_1899); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1901 = 7'h4f == data1Frac_14 ? $signed(8'sh2a) : $signed(_GEN_1900); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1902 = 7'h50 == data1Frac_14 ? $signed(8'sh29) : $signed(_GEN_1901); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1903 = 7'h51 == data1Frac_14 ? $signed(8'sh29) : $signed(_GEN_1902); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1904 = 7'h52 == data1Frac_14 ? $signed(8'sh29) : $signed(_GEN_1903); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1905 = 7'h53 == data1Frac_14 ? $signed(8'sh29) : $signed(_GEN_1904); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1906 = 7'h54 == data1Frac_14 ? $signed(8'sh29) : $signed(_GEN_1905); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1907 = 7'h55 == data1Frac_14 ? $signed(8'sh28) : $signed(_GEN_1906); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1908 = 7'h56 == data1Frac_14 ? $signed(8'sh28) : $signed(_GEN_1907); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1909 = 7'h57 == data1Frac_14 ? $signed(8'sh28) : $signed(_GEN_1908); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1910 = 7'h58 == data1Frac_14 ? $signed(8'sh28) : $signed(_GEN_1909); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1911 = 7'h59 == data1Frac_14 ? $signed(8'sh28) : $signed(_GEN_1910); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1912 = 7'h5a == data1Frac_14 ? $signed(8'sh27) : $signed(_GEN_1911); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1913 = 7'h5b == data1Frac_14 ? $signed(8'sh27) : $signed(_GEN_1912); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1914 = 7'h5c == data1Frac_14 ? $signed(8'sh27) : $signed(_GEN_1913); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1915 = 7'h5d == data1Frac_14 ? $signed(8'sh27) : $signed(_GEN_1914); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1916 = 7'h5e == data1Frac_14 ? $signed(8'sh26) : $signed(_GEN_1915); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1917 = 7'h5f == data1Frac_14 ? $signed(8'sh26) : $signed(_GEN_1916); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1918 = 7'h60 == data1Frac_14 ? $signed(8'sh26) : $signed(_GEN_1917); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1919 = 7'h61 == data1Frac_14 ? $signed(8'sh26) : $signed(_GEN_1918); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1920 = 7'h62 == data1Frac_14 ? $signed(8'sh26) : $signed(_GEN_1919); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1921 = 7'h63 == data1Frac_14 ? $signed(8'sh25) : $signed(_GEN_1920); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1922 = 7'h64 == data1Frac_14 ? $signed(8'sh25) : $signed(_GEN_1921); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1923 = 7'h65 == data1Frac_14 ? $signed(8'sh25) : $signed(_GEN_1922); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1924 = 7'h66 == data1Frac_14 ? $signed(8'sh25) : $signed(_GEN_1923); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1925 = 7'h67 == data1Frac_14 ? $signed(8'sh25) : $signed(_GEN_1924); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1926 = 7'h68 == data1Frac_14 ? $signed(8'sh24) : $signed(_GEN_1925); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1927 = 7'h69 == data1Frac_14 ? $signed(8'sh24) : $signed(_GEN_1926); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1928 = 7'h6a == data1Frac_14 ? $signed(8'sh24) : $signed(_GEN_1927); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1929 = 7'h6b == data1Frac_14 ? $signed(8'sh24) : $signed(_GEN_1928); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1930 = 7'h6c == data1Frac_14 ? $signed(8'sh24) : $signed(_GEN_1929); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1931 = 7'h6d == data1Frac_14 ? $signed(8'sh23) : $signed(_GEN_1930); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1932 = 7'h6e == data1Frac_14 ? $signed(8'sh23) : $signed(_GEN_1931); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1933 = 7'h6f == data1Frac_14 ? $signed(8'sh23) : $signed(_GEN_1932); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1934 = 7'h70 == data1Frac_14 ? $signed(8'sh23) : $signed(_GEN_1933); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1935 = 7'h71 == data1Frac_14 ? $signed(8'sh23) : $signed(_GEN_1934); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1936 = 7'h72 == data1Frac_14 ? $signed(8'sh23) : $signed(_GEN_1935); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1937 = 7'h73 == data1Frac_14 ? $signed(8'sh22) : $signed(_GEN_1936); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1938 = 7'h74 == data1Frac_14 ? $signed(8'sh22) : $signed(_GEN_1937); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1939 = 7'h75 == data1Frac_14 ? $signed(8'sh22) : $signed(_GEN_1938); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1940 = 7'h76 == data1Frac_14 ? $signed(8'sh22) : $signed(_GEN_1939); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1941 = 7'h77 == data1Frac_14 ? $signed(8'sh22) : $signed(_GEN_1940); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1942 = 7'h78 == data1Frac_14 ? $signed(8'sh21) : $signed(_GEN_1941); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1943 = 7'h79 == data1Frac_14 ? $signed(8'sh21) : $signed(_GEN_1942); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1944 = 7'h7a == data1Frac_14 ? $signed(8'sh21) : $signed(_GEN_1943); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1945 = 7'h7b == data1Frac_14 ? $signed(8'sh21) : $signed(_GEN_1944); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1946 = 7'h7c == data1Frac_14 ? $signed(8'sh21) : $signed(_GEN_1945); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1947 = 7'h7d == data1Frac_14 ? $signed(8'sh21) : $signed(_GEN_1946); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1948 = 7'h7e == data1Frac_14 ? $signed(8'sh20) : $signed(_GEN_1947); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1949 = 7'h7f == data1Frac_14 ? $signed(8'sh20) : $signed(_GEN_1948); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_44 = $signed(_GEN_1949) >>> data1Int_14; // @[exponent.scala 38:85]
  reg [7:0] data2_14; // @[Reg.scala 16:16]
  wire [7:0] _GEN_1953 = 7'h2 == data1Frac_15 ? $signed(8'sh3f) : $signed(8'sh40); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1954 = 7'h3 == data1Frac_15 ? $signed(8'sh3f) : $signed(_GEN_1953); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1955 = 7'h4 == data1Frac_15 ? $signed(8'sh3f) : $signed(_GEN_1954); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1956 = 7'h5 == data1Frac_15 ? $signed(8'sh3e) : $signed(_GEN_1955); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1957 = 7'h6 == data1Frac_15 ? $signed(8'sh3e) : $signed(_GEN_1956); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1958 = 7'h7 == data1Frac_15 ? $signed(8'sh3e) : $signed(_GEN_1957); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1959 = 7'h8 == data1Frac_15 ? $signed(8'sh3d) : $signed(_GEN_1958); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1960 = 7'h9 == data1Frac_15 ? $signed(8'sh3d) : $signed(_GEN_1959); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1961 = 7'ha == data1Frac_15 ? $signed(8'sh3d) : $signed(_GEN_1960); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1962 = 7'hb == data1Frac_15 ? $signed(8'sh3c) : $signed(_GEN_1961); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1963 = 7'hc == data1Frac_15 ? $signed(8'sh3c) : $signed(_GEN_1962); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1964 = 7'hd == data1Frac_15 ? $signed(8'sh3c) : $signed(_GEN_1963); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1965 = 7'he == data1Frac_15 ? $signed(8'sh3b) : $signed(_GEN_1964); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1966 = 7'hf == data1Frac_15 ? $signed(8'sh3b) : $signed(_GEN_1965); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1967 = 7'h10 == data1Frac_15 ? $signed(8'sh3b) : $signed(_GEN_1966); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1968 = 7'h11 == data1Frac_15 ? $signed(8'sh3a) : $signed(_GEN_1967); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1969 = 7'h12 == data1Frac_15 ? $signed(8'sh3a) : $signed(_GEN_1968); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1970 = 7'h13 == data1Frac_15 ? $signed(8'sh3a) : $signed(_GEN_1969); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1971 = 7'h14 == data1Frac_15 ? $signed(8'sh39) : $signed(_GEN_1970); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1972 = 7'h15 == data1Frac_15 ? $signed(8'sh39) : $signed(_GEN_1971); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1973 = 7'h16 == data1Frac_15 ? $signed(8'sh39) : $signed(_GEN_1972); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1974 = 7'h17 == data1Frac_15 ? $signed(8'sh39) : $signed(_GEN_1973); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1975 = 7'h18 == data1Frac_15 ? $signed(8'sh38) : $signed(_GEN_1974); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1976 = 7'h19 == data1Frac_15 ? $signed(8'sh38) : $signed(_GEN_1975); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1977 = 7'h1a == data1Frac_15 ? $signed(8'sh38) : $signed(_GEN_1976); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1978 = 7'h1b == data1Frac_15 ? $signed(8'sh37) : $signed(_GEN_1977); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1979 = 7'h1c == data1Frac_15 ? $signed(8'sh37) : $signed(_GEN_1978); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1980 = 7'h1d == data1Frac_15 ? $signed(8'sh37) : $signed(_GEN_1979); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1981 = 7'h1e == data1Frac_15 ? $signed(8'sh36) : $signed(_GEN_1980); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1982 = 7'h1f == data1Frac_15 ? $signed(8'sh36) : $signed(_GEN_1981); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1983 = 7'h20 == data1Frac_15 ? $signed(8'sh36) : $signed(_GEN_1982); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1984 = 7'h21 == data1Frac_15 ? $signed(8'sh36) : $signed(_GEN_1983); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1985 = 7'h22 == data1Frac_15 ? $signed(8'sh35) : $signed(_GEN_1984); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1986 = 7'h23 == data1Frac_15 ? $signed(8'sh35) : $signed(_GEN_1985); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1987 = 7'h24 == data1Frac_15 ? $signed(8'sh35) : $signed(_GEN_1986); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1988 = 7'h25 == data1Frac_15 ? $signed(8'sh34) : $signed(_GEN_1987); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1989 = 7'h26 == data1Frac_15 ? $signed(8'sh34) : $signed(_GEN_1988); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1990 = 7'h27 == data1Frac_15 ? $signed(8'sh34) : $signed(_GEN_1989); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1991 = 7'h28 == data1Frac_15 ? $signed(8'sh34) : $signed(_GEN_1990); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1992 = 7'h29 == data1Frac_15 ? $signed(8'sh33) : $signed(_GEN_1991); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1993 = 7'h2a == data1Frac_15 ? $signed(8'sh33) : $signed(_GEN_1992); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1994 = 7'h2b == data1Frac_15 ? $signed(8'sh33) : $signed(_GEN_1993); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1995 = 7'h2c == data1Frac_15 ? $signed(8'sh32) : $signed(_GEN_1994); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1996 = 7'h2d == data1Frac_15 ? $signed(8'sh32) : $signed(_GEN_1995); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1997 = 7'h2e == data1Frac_15 ? $signed(8'sh32) : $signed(_GEN_1996); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1998 = 7'h2f == data1Frac_15 ? $signed(8'sh32) : $signed(_GEN_1997); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_1999 = 7'h30 == data1Frac_15 ? $signed(8'sh31) : $signed(_GEN_1998); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2000 = 7'h31 == data1Frac_15 ? $signed(8'sh31) : $signed(_GEN_1999); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2001 = 7'h32 == data1Frac_15 ? $signed(8'sh31) : $signed(_GEN_2000); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2002 = 7'h33 == data1Frac_15 ? $signed(8'sh31) : $signed(_GEN_2001); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2003 = 7'h34 == data1Frac_15 ? $signed(8'sh30) : $signed(_GEN_2002); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2004 = 7'h35 == data1Frac_15 ? $signed(8'sh30) : $signed(_GEN_2003); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2005 = 7'h36 == data1Frac_15 ? $signed(8'sh30) : $signed(_GEN_2004); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2006 = 7'h37 == data1Frac_15 ? $signed(8'sh30) : $signed(_GEN_2005); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2007 = 7'h38 == data1Frac_15 ? $signed(8'sh2f) : $signed(_GEN_2006); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2008 = 7'h39 == data1Frac_15 ? $signed(8'sh2f) : $signed(_GEN_2007); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2009 = 7'h3a == data1Frac_15 ? $signed(8'sh2f) : $signed(_GEN_2008); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2010 = 7'h3b == data1Frac_15 ? $signed(8'sh2e) : $signed(_GEN_2009); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2011 = 7'h3c == data1Frac_15 ? $signed(8'sh2e) : $signed(_GEN_2010); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2012 = 7'h3d == data1Frac_15 ? $signed(8'sh2e) : $signed(_GEN_2011); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2013 = 7'h3e == data1Frac_15 ? $signed(8'sh2e) : $signed(_GEN_2012); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2014 = 7'h3f == data1Frac_15 ? $signed(8'sh2e) : $signed(_GEN_2013); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2015 = 7'h40 == data1Frac_15 ? $signed(8'sh2d) : $signed(_GEN_2014); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2016 = 7'h41 == data1Frac_15 ? $signed(8'sh2d) : $signed(_GEN_2015); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2017 = 7'h42 == data1Frac_15 ? $signed(8'sh2d) : $signed(_GEN_2016); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2018 = 7'h43 == data1Frac_15 ? $signed(8'sh2d) : $signed(_GEN_2017); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2019 = 7'h44 == data1Frac_15 ? $signed(8'sh2c) : $signed(_GEN_2018); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2020 = 7'h45 == data1Frac_15 ? $signed(8'sh2c) : $signed(_GEN_2019); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2021 = 7'h46 == data1Frac_15 ? $signed(8'sh2c) : $signed(_GEN_2020); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2022 = 7'h47 == data1Frac_15 ? $signed(8'sh2c) : $signed(_GEN_2021); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2023 = 7'h48 == data1Frac_15 ? $signed(8'sh2b) : $signed(_GEN_2022); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2024 = 7'h49 == data1Frac_15 ? $signed(8'sh2b) : $signed(_GEN_2023); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2025 = 7'h4a == data1Frac_15 ? $signed(8'sh2b) : $signed(_GEN_2024); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2026 = 7'h4b == data1Frac_15 ? $signed(8'sh2b) : $signed(_GEN_2025); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2027 = 7'h4c == data1Frac_15 ? $signed(8'sh2a) : $signed(_GEN_2026); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2028 = 7'h4d == data1Frac_15 ? $signed(8'sh2a) : $signed(_GEN_2027); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2029 = 7'h4e == data1Frac_15 ? $signed(8'sh2a) : $signed(_GEN_2028); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2030 = 7'h4f == data1Frac_15 ? $signed(8'sh2a) : $signed(_GEN_2029); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2031 = 7'h50 == data1Frac_15 ? $signed(8'sh29) : $signed(_GEN_2030); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2032 = 7'h51 == data1Frac_15 ? $signed(8'sh29) : $signed(_GEN_2031); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2033 = 7'h52 == data1Frac_15 ? $signed(8'sh29) : $signed(_GEN_2032); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2034 = 7'h53 == data1Frac_15 ? $signed(8'sh29) : $signed(_GEN_2033); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2035 = 7'h54 == data1Frac_15 ? $signed(8'sh29) : $signed(_GEN_2034); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2036 = 7'h55 == data1Frac_15 ? $signed(8'sh28) : $signed(_GEN_2035); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2037 = 7'h56 == data1Frac_15 ? $signed(8'sh28) : $signed(_GEN_2036); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2038 = 7'h57 == data1Frac_15 ? $signed(8'sh28) : $signed(_GEN_2037); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2039 = 7'h58 == data1Frac_15 ? $signed(8'sh28) : $signed(_GEN_2038); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2040 = 7'h59 == data1Frac_15 ? $signed(8'sh28) : $signed(_GEN_2039); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2041 = 7'h5a == data1Frac_15 ? $signed(8'sh27) : $signed(_GEN_2040); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2042 = 7'h5b == data1Frac_15 ? $signed(8'sh27) : $signed(_GEN_2041); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2043 = 7'h5c == data1Frac_15 ? $signed(8'sh27) : $signed(_GEN_2042); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2044 = 7'h5d == data1Frac_15 ? $signed(8'sh27) : $signed(_GEN_2043); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2045 = 7'h5e == data1Frac_15 ? $signed(8'sh26) : $signed(_GEN_2044); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2046 = 7'h5f == data1Frac_15 ? $signed(8'sh26) : $signed(_GEN_2045); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2047 = 7'h60 == data1Frac_15 ? $signed(8'sh26) : $signed(_GEN_2046); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2048 = 7'h61 == data1Frac_15 ? $signed(8'sh26) : $signed(_GEN_2047); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2049 = 7'h62 == data1Frac_15 ? $signed(8'sh26) : $signed(_GEN_2048); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2050 = 7'h63 == data1Frac_15 ? $signed(8'sh25) : $signed(_GEN_2049); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2051 = 7'h64 == data1Frac_15 ? $signed(8'sh25) : $signed(_GEN_2050); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2052 = 7'h65 == data1Frac_15 ? $signed(8'sh25) : $signed(_GEN_2051); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2053 = 7'h66 == data1Frac_15 ? $signed(8'sh25) : $signed(_GEN_2052); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2054 = 7'h67 == data1Frac_15 ? $signed(8'sh25) : $signed(_GEN_2053); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2055 = 7'h68 == data1Frac_15 ? $signed(8'sh24) : $signed(_GEN_2054); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2056 = 7'h69 == data1Frac_15 ? $signed(8'sh24) : $signed(_GEN_2055); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2057 = 7'h6a == data1Frac_15 ? $signed(8'sh24) : $signed(_GEN_2056); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2058 = 7'h6b == data1Frac_15 ? $signed(8'sh24) : $signed(_GEN_2057); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2059 = 7'h6c == data1Frac_15 ? $signed(8'sh24) : $signed(_GEN_2058); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2060 = 7'h6d == data1Frac_15 ? $signed(8'sh23) : $signed(_GEN_2059); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2061 = 7'h6e == data1Frac_15 ? $signed(8'sh23) : $signed(_GEN_2060); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2062 = 7'h6f == data1Frac_15 ? $signed(8'sh23) : $signed(_GEN_2061); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2063 = 7'h70 == data1Frac_15 ? $signed(8'sh23) : $signed(_GEN_2062); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2064 = 7'h71 == data1Frac_15 ? $signed(8'sh23) : $signed(_GEN_2063); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2065 = 7'h72 == data1Frac_15 ? $signed(8'sh23) : $signed(_GEN_2064); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2066 = 7'h73 == data1Frac_15 ? $signed(8'sh22) : $signed(_GEN_2065); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2067 = 7'h74 == data1Frac_15 ? $signed(8'sh22) : $signed(_GEN_2066); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2068 = 7'h75 == data1Frac_15 ? $signed(8'sh22) : $signed(_GEN_2067); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2069 = 7'h76 == data1Frac_15 ? $signed(8'sh22) : $signed(_GEN_2068); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2070 = 7'h77 == data1Frac_15 ? $signed(8'sh22) : $signed(_GEN_2069); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2071 = 7'h78 == data1Frac_15 ? $signed(8'sh21) : $signed(_GEN_2070); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2072 = 7'h79 == data1Frac_15 ? $signed(8'sh21) : $signed(_GEN_2071); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2073 = 7'h7a == data1Frac_15 ? $signed(8'sh21) : $signed(_GEN_2072); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2074 = 7'h7b == data1Frac_15 ? $signed(8'sh21) : $signed(_GEN_2073); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2075 = 7'h7c == data1Frac_15 ? $signed(8'sh21) : $signed(_GEN_2074); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2076 = 7'h7d == data1Frac_15 ? $signed(8'sh21) : $signed(_GEN_2075); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2077 = 7'h7e == data1Frac_15 ? $signed(8'sh20) : $signed(_GEN_2076); // @[exponent.scala 38:{47,47}]
  wire [7:0] _GEN_2078 = 7'h7f == data1Frac_15 ? $signed(8'sh20) : $signed(_GEN_2077); // @[exponent.scala 38:{47,47}]
  wire [7:0] _data2_T_47 = $signed(_GEN_2078) >>> data1Int_15; // @[exponent.scala 38:85]
  reg [7:0] data2_15; // @[Reg.scala 16:16]
  PipelineHsk hsk ( // @[exponent.scala 20:21]
    .clock(hsk_clock),
    .reset(hsk_reset),
    .io_validPre(hsk_io_validPre),
    .io_readyPre(hsk_io_readyPre),
    .io_lastPre(hsk_io_lastPre),
    .io_validNxt(hsk_io_validNxt),
    .io_readyNxt(hsk_io_readyNxt),
    .io_regen_0(hsk_io_regen_0),
    .io_regen_1(hsk_io_regen_1),
    .io_lastNxt(hsk_io_lastNxt)
  );
  assign io_input_ready = hsk_io_readyPre; // @[exponent.scala 22:20]
  assign io_output_valid = hsk_io_validNxt; // @[exponent.scala 23:21]
  assign io_output_bits_x_0 = data2_0; // @[exponent.scala 40:22]
  assign io_output_bits_x_1 = data2_1; // @[exponent.scala 40:22]
  assign io_output_bits_x_2 = data2_2; // @[exponent.scala 40:22]
  assign io_output_bits_x_3 = data2_3; // @[exponent.scala 40:22]
  assign io_output_bits_x_4 = data2_4; // @[exponent.scala 40:22]
  assign io_output_bits_x_5 = data2_5; // @[exponent.scala 40:22]
  assign io_output_bits_x_6 = data2_6; // @[exponent.scala 40:22]
  assign io_output_bits_x_7 = data2_7; // @[exponent.scala 40:22]
  assign io_output_bits_x_8 = data2_8; // @[exponent.scala 40:22]
  assign io_output_bits_x_9 = data2_9; // @[exponent.scala 40:22]
  assign io_output_bits_x_10 = data2_10; // @[exponent.scala 40:22]
  assign io_output_bits_x_11 = data2_11; // @[exponent.scala 40:22]
  assign io_output_bits_x_12 = data2_12; // @[exponent.scala 40:22]
  assign io_output_bits_x_13 = data2_13; // @[exponent.scala 40:22]
  assign io_output_bits_x_14 = data2_14; // @[exponent.scala 40:22]
  assign io_output_bits_x_15 = data2_15; // @[exponent.scala 40:22]
  assign io_output_bits_last = hsk_io_lastNxt; // @[exponent.scala 26:25]
  assign hsk_clock = clock;
  assign hsk_reset = reset;
  assign hsk_io_validPre = io_input_valid; // @[exponent.scala 21:21]
  assign hsk_io_lastPre = io_input_bits_last; // @[exponent.scala 25:20]
  assign hsk_io_readyNxt = io_output_ready; // @[exponent.scala 24:21]
  always @(posedge clock) begin
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_0 <= _data1_T; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_1 <= _data1_T_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_2 <= _data1_T_2; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_3 <= _data1_T_3; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_4 <= _data1_T_4; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_5 <= _data1_T_5; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_6 <= _data1_T_6; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_7 <= _data1_T_7; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_8 <= _data1_T_8; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_9 <= _data1_T_9; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_10 <= _data1_T_10; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_11 <= _data1_T_11; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_12 <= _data1_T_12; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_13 <= _data1_T_13; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_14 <= _data1_T_14; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1_15 <= _data1_T_15; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_0 <= _data2_T_2; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_1 <= _data2_T_5; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_2 <= _data2_T_8; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_3 <= _data2_T_11; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_4 <= _data2_T_14; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_5 <= _data2_T_17; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_6 <= _data2_T_20; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_7 <= _data2_T_23; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_8 <= _data2_T_26; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_9 <= _data2_T_29; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_10 <= _data2_T_32; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_11 <= _data2_T_35; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_12 <= _data2_T_38; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_13 <= _data2_T_41; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_14 <= _data2_T_44; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2_15 <= _data2_T_47; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data1_0 = _RAND_0[12:0];
  _RAND_1 = {1{`RANDOM}};
  data1_1 = _RAND_1[12:0];
  _RAND_2 = {1{`RANDOM}};
  data1_2 = _RAND_2[12:0];
  _RAND_3 = {1{`RANDOM}};
  data1_3 = _RAND_3[12:0];
  _RAND_4 = {1{`RANDOM}};
  data1_4 = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  data1_5 = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  data1_6 = _RAND_6[12:0];
  _RAND_7 = {1{`RANDOM}};
  data1_7 = _RAND_7[12:0];
  _RAND_8 = {1{`RANDOM}};
  data1_8 = _RAND_8[12:0];
  _RAND_9 = {1{`RANDOM}};
  data1_9 = _RAND_9[12:0];
  _RAND_10 = {1{`RANDOM}};
  data1_10 = _RAND_10[12:0];
  _RAND_11 = {1{`RANDOM}};
  data1_11 = _RAND_11[12:0];
  _RAND_12 = {1{`RANDOM}};
  data1_12 = _RAND_12[12:0];
  _RAND_13 = {1{`RANDOM}};
  data1_13 = _RAND_13[12:0];
  _RAND_14 = {1{`RANDOM}};
  data1_14 = _RAND_14[12:0];
  _RAND_15 = {1{`RANDOM}};
  data1_15 = _RAND_15[12:0];
  _RAND_16 = {1{`RANDOM}};
  data2_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data2_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data2_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data2_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data2_4 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data2_5 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data2_6 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data2_7 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data2_8 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data2_9 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data2_10 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data2_11 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data2_12 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data2_13 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data2_14 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data2_15 = _RAND_31[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Hsk1ton(
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_0_x_0,
  input  [7:0] io_input_bits_0_x_1,
  input  [7:0] io_input_bits_0_x_2,
  input  [7:0] io_input_bits_0_x_3,
  input  [7:0] io_input_bits_0_x_4,
  input  [7:0] io_input_bits_0_x_5,
  input  [7:0] io_input_bits_0_x_6,
  input  [7:0] io_input_bits_0_x_7,
  input  [7:0] io_input_bits_0_x_8,
  input  [7:0] io_input_bits_0_x_9,
  input  [7:0] io_input_bits_0_x_10,
  input  [7:0] io_input_bits_0_x_11,
  input  [7:0] io_input_bits_0_x_12,
  input  [7:0] io_input_bits_0_x_13,
  input  [7:0] io_input_bits_0_x_14,
  input  [7:0] io_input_bits_0_x_15,
  input        io_input_bits_0_last,
  input  [7:0] io_input_bits_1_x_0,
  input  [7:0] io_input_bits_1_x_1,
  input  [7:0] io_input_bits_1_x_2,
  input  [7:0] io_input_bits_1_x_3,
  input  [7:0] io_input_bits_1_x_4,
  input  [7:0] io_input_bits_1_x_5,
  input  [7:0] io_input_bits_1_x_6,
  input  [7:0] io_input_bits_1_x_7,
  input  [7:0] io_input_bits_1_x_8,
  input  [7:0] io_input_bits_1_x_9,
  input  [7:0] io_input_bits_1_x_10,
  input  [7:0] io_input_bits_1_x_11,
  input  [7:0] io_input_bits_1_x_12,
  input  [7:0] io_input_bits_1_x_13,
  input  [7:0] io_input_bits_1_x_14,
  input  [7:0] io_input_bits_1_x_15,
  input        io_input_bits_1_last,
  input        io_output_0_ready,
  output       io_output_0_valid,
  output [7:0] io_output_0_bits_x_0,
  output [7:0] io_output_0_bits_x_1,
  output [7:0] io_output_0_bits_x_2,
  output [7:0] io_output_0_bits_x_3,
  output [7:0] io_output_0_bits_x_4,
  output [7:0] io_output_0_bits_x_5,
  output [7:0] io_output_0_bits_x_6,
  output [7:0] io_output_0_bits_x_7,
  output [7:0] io_output_0_bits_x_8,
  output [7:0] io_output_0_bits_x_9,
  output [7:0] io_output_0_bits_x_10,
  output [7:0] io_output_0_bits_x_11,
  output [7:0] io_output_0_bits_x_12,
  output [7:0] io_output_0_bits_x_13,
  output [7:0] io_output_0_bits_x_14,
  output [7:0] io_output_0_bits_x_15,
  output       io_output_0_bits_last,
  input        io_output_1_ready,
  output       io_output_1_valid,
  output [7:0] io_output_1_bits_x_0,
  output [7:0] io_output_1_bits_x_1,
  output [7:0] io_output_1_bits_x_2,
  output [7:0] io_output_1_bits_x_3,
  output [7:0] io_output_1_bits_x_4,
  output [7:0] io_output_1_bits_x_5,
  output [7:0] io_output_1_bits_x_6,
  output [7:0] io_output_1_bits_x_7,
  output [7:0] io_output_1_bits_x_8,
  output [7:0] io_output_1_bits_x_9,
  output [7:0] io_output_1_bits_x_10,
  output [7:0] io_output_1_bits_x_11,
  output [7:0] io_output_1_bits_x_12,
  output [7:0] io_output_1_bits_x_13,
  output [7:0] io_output_1_bits_x_14,
  output [7:0] io_output_1_bits_x_15,
  output       io_output_1_bits_last
);
  assign io_input_ready = io_output_0_ready & io_output_1_ready; // @[hsk1ton.scala 12:58]
  assign io_output_0_valid = io_input_valid & (~io_output_0_ready | io_output_1_ready); // @[hsk1ton.scala 14:72]
  assign io_output_0_bits_x_0 = io_input_bits_0_x_0; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_1 = io_input_bits_0_x_1; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_2 = io_input_bits_0_x_2; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_3 = io_input_bits_0_x_3; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_4 = io_input_bits_0_x_4; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_5 = io_input_bits_0_x_5; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_6 = io_input_bits_0_x_6; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_7 = io_input_bits_0_x_7; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_8 = io_input_bits_0_x_8; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_9 = io_input_bits_0_x_9; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_10 = io_input_bits_0_x_10; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_11 = io_input_bits_0_x_11; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_12 = io_input_bits_0_x_12; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_13 = io_input_bits_0_x_13; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_14 = io_input_bits_0_x_14; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_15 = io_input_bits_0_x_15; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_last = io_input_bits_0_last; // @[hsk1ton.scala 13:54]
  assign io_output_1_valid = io_input_valid & (~io_output_1_ready | io_output_0_ready); // @[hsk1ton.scala 14:72]
  assign io_output_1_bits_x_0 = io_input_bits_1_x_0; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_1 = io_input_bits_1_x_1; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_2 = io_input_bits_1_x_2; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_3 = io_input_bits_1_x_3; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_4 = io_input_bits_1_x_4; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_5 = io_input_bits_1_x_5; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_6 = io_input_bits_1_x_6; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_7 = io_input_bits_1_x_7; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_8 = io_input_bits_1_x_8; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_9 = io_input_bits_1_x_9; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_10 = io_input_bits_1_x_10; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_11 = io_input_bits_1_x_11; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_12 = io_input_bits_1_x_12; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_13 = io_input_bits_1_x_13; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_14 = io_input_bits_1_x_14; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_15 = io_input_bits_1_x_15; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_last = io_input_bits_1_last; // @[hsk1ton.scala 13:54]
endmodule
module Arbiternto1(
  output       io_input_0_ready,
  input        io_input_0_valid,
  input  [7:0] io_input_0_bits_x_0,
  input  [7:0] io_input_0_bits_x_1,
  input  [7:0] io_input_0_bits_x_2,
  input  [7:0] io_input_0_bits_x_3,
  input  [7:0] io_input_0_bits_x_4,
  input  [7:0] io_input_0_bits_x_5,
  input  [7:0] io_input_0_bits_x_6,
  input  [7:0] io_input_0_bits_x_7,
  input  [7:0] io_input_0_bits_x_8,
  input  [7:0] io_input_0_bits_x_9,
  input  [7:0] io_input_0_bits_x_10,
  input  [7:0] io_input_0_bits_x_11,
  input  [7:0] io_input_0_bits_x_12,
  input  [7:0] io_input_0_bits_x_13,
  input  [7:0] io_input_0_bits_x_14,
  input  [7:0] io_input_0_bits_x_15,
  input        io_input_0_bits_last,
  output       io_input_1_ready,
  input        io_input_1_valid,
  input  [7:0] io_input_1_bits_x_0,
  input  [7:0] io_input_1_bits_x_1,
  input  [7:0] io_input_1_bits_x_2,
  input  [7:0] io_input_1_bits_x_3,
  input  [7:0] io_input_1_bits_x_4,
  input  [7:0] io_input_1_bits_x_5,
  input  [7:0] io_input_1_bits_x_6,
  input  [7:0] io_input_1_bits_x_7,
  input  [7:0] io_input_1_bits_x_8,
  input  [7:0] io_input_1_bits_x_9,
  input  [7:0] io_input_1_bits_x_10,
  input  [7:0] io_input_1_bits_x_11,
  input  [7:0] io_input_1_bits_x_12,
  input  [7:0] io_input_1_bits_x_13,
  input  [7:0] io_input_1_bits_x_14,
  input  [7:0] io_input_1_bits_x_15,
  input        io_input_1_bits_last,
  input        io_sel,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_x_0,
  output [7:0] io_output_bits_x_1,
  output [7:0] io_output_bits_x_2,
  output [7:0] io_output_bits_x_3,
  output [7:0] io_output_bits_x_4,
  output [7:0] io_output_bits_x_5,
  output [7:0] io_output_bits_x_6,
  output [7:0] io_output_bits_x_7,
  output [7:0] io_output_bits_x_8,
  output [7:0] io_output_bits_x_9,
  output [7:0] io_output_bits_x_10,
  output [7:0] io_output_bits_x_11,
  output [7:0] io_output_bits_x_12,
  output [7:0] io_output_bits_x_13,
  output [7:0] io_output_bits_x_14,
  output [7:0] io_output_bits_x_15,
  output       io_output_bits_last
);
  assign io_input_0_ready = ~io_sel & io_output_ready; // @[arbiternto1.scala 17:44]
  assign io_input_1_ready = io_sel & io_output_ready; // @[arbiternto1.scala 17:44]
  assign io_output_valid = io_sel ? io_input_1_valid : io_input_0_valid; // @[arbiternto1.scala 15:{21,21}]
  assign io_output_bits_x_0 = io_sel ? $signed(io_input_1_bits_x_0) : $signed(io_input_0_bits_x_0); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_1 = io_sel ? $signed(io_input_1_bits_x_1) : $signed(io_input_0_bits_x_1); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_2 = io_sel ? $signed(io_input_1_bits_x_2) : $signed(io_input_0_bits_x_2); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_3 = io_sel ? $signed(io_input_1_bits_x_3) : $signed(io_input_0_bits_x_3); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_4 = io_sel ? $signed(io_input_1_bits_x_4) : $signed(io_input_0_bits_x_4); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_5 = io_sel ? $signed(io_input_1_bits_x_5) : $signed(io_input_0_bits_x_5); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_6 = io_sel ? $signed(io_input_1_bits_x_6) : $signed(io_input_0_bits_x_6); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_7 = io_sel ? $signed(io_input_1_bits_x_7) : $signed(io_input_0_bits_x_7); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_8 = io_sel ? $signed(io_input_1_bits_x_8) : $signed(io_input_0_bits_x_8); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_9 = io_sel ? $signed(io_input_1_bits_x_9) : $signed(io_input_0_bits_x_9); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_10 = io_sel ? $signed(io_input_1_bits_x_10) : $signed(io_input_0_bits_x_10); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_11 = io_sel ? $signed(io_input_1_bits_x_11) : $signed(io_input_0_bits_x_11); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_12 = io_sel ? $signed(io_input_1_bits_x_12) : $signed(io_input_0_bits_x_12); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_13 = io_sel ? $signed(io_input_1_bits_x_13) : $signed(io_input_0_bits_x_13); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_14 = io_sel ? $signed(io_input_1_bits_x_14) : $signed(io_input_0_bits_x_14); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_x_15 = io_sel ? $signed(io_input_1_bits_x_15) : $signed(io_input_0_bits_x_15); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_last = io_sel ? io_input_1_bits_last : io_input_0_bits_last; // @[arbiternto1.scala 14:{20,20}]
endmodule
module Arbiter1ton(
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_x_0,
  input  [7:0] io_input_bits_x_1,
  input  [7:0] io_input_bits_x_2,
  input  [7:0] io_input_bits_x_3,
  input  [7:0] io_input_bits_x_4,
  input  [7:0] io_input_bits_x_5,
  input  [7:0] io_input_bits_x_6,
  input  [7:0] io_input_bits_x_7,
  input  [7:0] io_input_bits_x_8,
  input  [7:0] io_input_bits_x_9,
  input  [7:0] io_input_bits_x_10,
  input  [7:0] io_input_bits_x_11,
  input  [7:0] io_input_bits_x_12,
  input  [7:0] io_input_bits_x_13,
  input  [7:0] io_input_bits_x_14,
  input  [7:0] io_input_bits_x_15,
  input        io_input_bits_last,
  input        io_sel,
  input        io_output_0_ready,
  output       io_output_0_valid,
  output [7:0] io_output_0_bits_x_0,
  output [7:0] io_output_0_bits_x_1,
  output [7:0] io_output_0_bits_x_2,
  output [7:0] io_output_0_bits_x_3,
  output [7:0] io_output_0_bits_x_4,
  output [7:0] io_output_0_bits_x_5,
  output [7:0] io_output_0_bits_x_6,
  output [7:0] io_output_0_bits_x_7,
  output [7:0] io_output_0_bits_x_8,
  output [7:0] io_output_0_bits_x_9,
  output [7:0] io_output_0_bits_x_10,
  output [7:0] io_output_0_bits_x_11,
  output [7:0] io_output_0_bits_x_12,
  output [7:0] io_output_0_bits_x_13,
  output [7:0] io_output_0_bits_x_14,
  output [7:0] io_output_0_bits_x_15,
  output       io_output_0_bits_last,
  input        io_output_1_ready,
  output       io_output_1_valid,
  output [7:0] io_output_1_bits_x_0,
  output [7:0] io_output_1_bits_x_1,
  output [7:0] io_output_1_bits_x_2,
  output [7:0] io_output_1_bits_x_3,
  output [7:0] io_output_1_bits_x_4,
  output [7:0] io_output_1_bits_x_5,
  output [7:0] io_output_1_bits_x_6,
  output [7:0] io_output_1_bits_x_7,
  output [7:0] io_output_1_bits_x_8,
  output [7:0] io_output_1_bits_x_9,
  output [7:0] io_output_1_bits_x_10,
  output [7:0] io_output_1_bits_x_11,
  output [7:0] io_output_1_bits_x_12,
  output [7:0] io_output_1_bits_x_13,
  output [7:0] io_output_1_bits_x_14,
  output [7:0] io_output_1_bits_x_15,
  output       io_output_1_bits_last
);
  assign io_input_ready = io_sel ? io_output_1_ready : io_output_0_ready; // @[arbiter1ton.scala 16:{20,20}]
  assign io_output_0_valid = ~io_sel & io_input_valid; // @[arbiter1ton.scala 18:44]
  assign io_output_0_bits_x_0 = io_input_bits_x_0; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_1 = io_input_bits_x_1; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_2 = io_input_bits_x_2; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_3 = io_input_bits_x_3; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_4 = io_input_bits_x_4; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_5 = io_input_bits_x_5; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_6 = io_input_bits_x_6; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_7 = io_input_bits_x_7; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_8 = io_input_bits_x_8; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_9 = io_input_bits_x_9; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_10 = io_input_bits_x_10; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_11 = io_input_bits_x_11; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_12 = io_input_bits_x_12; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_13 = io_input_bits_x_13; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_14 = io_input_bits_x_14; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_15 = io_input_bits_x_15; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_last = io_input_bits_last; // @[arbiter1ton.scala 19:26]
  assign io_output_1_valid = io_sel & io_input_valid; // @[arbiter1ton.scala 18:44]
  assign io_output_1_bits_x_0 = io_input_bits_x_0; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_1 = io_input_bits_x_1; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_2 = io_input_bits_x_2; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_3 = io_input_bits_x_3; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_4 = io_input_bits_x_4; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_5 = io_input_bits_x_5; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_6 = io_input_bits_x_6; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_7 = io_input_bits_x_7; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_8 = io_input_bits_x_8; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_9 = io_input_bits_x_9; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_10 = io_input_bits_x_10; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_11 = io_input_bits_x_11; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_12 = io_input_bits_x_12; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_13 = io_input_bits_x_13; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_14 = io_input_bits_x_14; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_x_15 = io_input_bits_x_15; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_last = io_input_bits_last; // @[arbiter1ton.scala 19:26]
endmodule
module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_x_0,
  input  [7:0] io_enq_bits_x_1,
  input  [7:0] io_enq_bits_x_2,
  input  [7:0] io_enq_bits_x_3,
  input  [7:0] io_enq_bits_x_4,
  input  [7:0] io_enq_bits_x_5,
  input  [7:0] io_enq_bits_x_6,
  input  [7:0] io_enq_bits_x_7,
  input  [7:0] io_enq_bits_x_8,
  input  [7:0] io_enq_bits_x_9,
  input  [7:0] io_enq_bits_x_10,
  input  [7:0] io_enq_bits_x_11,
  input  [7:0] io_enq_bits_x_12,
  input  [7:0] io_enq_bits_x_13,
  input  [7:0] io_enq_bits_x_14,
  input  [7:0] io_enq_bits_x_15,
  input        io_enq_bits_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_x_0,
  output [7:0] io_deq_bits_x_1,
  output [7:0] io_deq_bits_x_2,
  output [7:0] io_deq_bits_x_3,
  output [7:0] io_deq_bits_x_4,
  output [7:0] io_deq_bits_x_5,
  output [7:0] io_deq_bits_x_6,
  output [7:0] io_deq_bits_x_7,
  output [7:0] io_deq_bits_x_8,
  output [7:0] io_deq_bits_x_9,
  output [7:0] io_deq_bits_x_10,
  output [7:0] io_deq_bits_x_11,
  output [7:0] io_deq_bits_x_12,
  output [7:0] io_deq_bits_x_13,
  output [7:0] io_deq_bits_x_14,
  output [7:0] io_deq_bits_x_15,
  output       io_deq_bits_last
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_x_0 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_0_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_0_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_0_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_0_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_0_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_0_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_1 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_1_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_1_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_1_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_1_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_1_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_1_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_2 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_2_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_2_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_2_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_2_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_2_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_2_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_3 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_3_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_3_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_3_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_3_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_3_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_3_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_4 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_4_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_4_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_4_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_4_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_4_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_4_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_5 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_5_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_5_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_5_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_5_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_5_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_5_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_6 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_6_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_6_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_6_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_6_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_6_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_6_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_7 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_7_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_7_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_7_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_7_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_7_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_7_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_8 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_8_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_8_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_8_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_8_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_8_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_8_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_9 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_9_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_9_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_9_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_9_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_9_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_9_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_10 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_10_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_10_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_10_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_10_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_10_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_10_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_11 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_11_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_11_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_11_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_11_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_11_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_11_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_12 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_12_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_12_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_12_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_12_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_12_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_12_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_13 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_13_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_13_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_13_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_13_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_13_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_13_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_14 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_14_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_14_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_14_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_14_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_14_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_14_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_x_15 [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_x_15_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_x_15_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_x_15_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_x_15_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_x_15_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_x_15_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_x_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_0_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_0_io_deq_bits_MPORT_data = ram_x_0[ram_x_0_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_0_MPORT_data = io_enq_bits_x_0;
  assign ram_x_0_MPORT_addr = 1'h0;
  assign ram_x_0_MPORT_mask = 1'h1;
  assign ram_x_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_1_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_1_io_deq_bits_MPORT_data = ram_x_1[ram_x_1_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_1_MPORT_data = io_enq_bits_x_1;
  assign ram_x_1_MPORT_addr = 1'h0;
  assign ram_x_1_MPORT_mask = 1'h1;
  assign ram_x_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_2_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_2_io_deq_bits_MPORT_data = ram_x_2[ram_x_2_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_2_MPORT_data = io_enq_bits_x_2;
  assign ram_x_2_MPORT_addr = 1'h0;
  assign ram_x_2_MPORT_mask = 1'h1;
  assign ram_x_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_3_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_3_io_deq_bits_MPORT_data = ram_x_3[ram_x_3_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_3_MPORT_data = io_enq_bits_x_3;
  assign ram_x_3_MPORT_addr = 1'h0;
  assign ram_x_3_MPORT_mask = 1'h1;
  assign ram_x_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_4_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_4_io_deq_bits_MPORT_data = ram_x_4[ram_x_4_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_4_MPORT_data = io_enq_bits_x_4;
  assign ram_x_4_MPORT_addr = 1'h0;
  assign ram_x_4_MPORT_mask = 1'h1;
  assign ram_x_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_5_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_5_io_deq_bits_MPORT_data = ram_x_5[ram_x_5_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_5_MPORT_data = io_enq_bits_x_5;
  assign ram_x_5_MPORT_addr = 1'h0;
  assign ram_x_5_MPORT_mask = 1'h1;
  assign ram_x_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_6_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_6_io_deq_bits_MPORT_data = ram_x_6[ram_x_6_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_6_MPORT_data = io_enq_bits_x_6;
  assign ram_x_6_MPORT_addr = 1'h0;
  assign ram_x_6_MPORT_mask = 1'h1;
  assign ram_x_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_7_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_7_io_deq_bits_MPORT_data = ram_x_7[ram_x_7_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_7_MPORT_data = io_enq_bits_x_7;
  assign ram_x_7_MPORT_addr = 1'h0;
  assign ram_x_7_MPORT_mask = 1'h1;
  assign ram_x_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_8_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_8_io_deq_bits_MPORT_data = ram_x_8[ram_x_8_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_8_MPORT_data = io_enq_bits_x_8;
  assign ram_x_8_MPORT_addr = 1'h0;
  assign ram_x_8_MPORT_mask = 1'h1;
  assign ram_x_8_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_9_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_9_io_deq_bits_MPORT_data = ram_x_9[ram_x_9_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_9_MPORT_data = io_enq_bits_x_9;
  assign ram_x_9_MPORT_addr = 1'h0;
  assign ram_x_9_MPORT_mask = 1'h1;
  assign ram_x_9_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_10_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_10_io_deq_bits_MPORT_data = ram_x_10[ram_x_10_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_10_MPORT_data = io_enq_bits_x_10;
  assign ram_x_10_MPORT_addr = 1'h0;
  assign ram_x_10_MPORT_mask = 1'h1;
  assign ram_x_10_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_11_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_11_io_deq_bits_MPORT_data = ram_x_11[ram_x_11_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_11_MPORT_data = io_enq_bits_x_11;
  assign ram_x_11_MPORT_addr = 1'h0;
  assign ram_x_11_MPORT_mask = 1'h1;
  assign ram_x_11_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_12_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_12_io_deq_bits_MPORT_data = ram_x_12[ram_x_12_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_12_MPORT_data = io_enq_bits_x_12;
  assign ram_x_12_MPORT_addr = 1'h0;
  assign ram_x_12_MPORT_mask = 1'h1;
  assign ram_x_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_13_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_13_io_deq_bits_MPORT_data = ram_x_13[ram_x_13_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_13_MPORT_data = io_enq_bits_x_13;
  assign ram_x_13_MPORT_addr = 1'h0;
  assign ram_x_13_MPORT_mask = 1'h1;
  assign ram_x_13_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_14_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_14_io_deq_bits_MPORT_data = ram_x_14[ram_x_14_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_14_MPORT_data = io_enq_bits_x_14;
  assign ram_x_14_MPORT_addr = 1'h0;
  assign ram_x_14_MPORT_mask = 1'h1;
  assign ram_x_14_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_x_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_x_15_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_x_15_io_deq_bits_MPORT_data = ram_x_15[ram_x_15_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_x_15_MPORT_data = io_enq_bits_x_15;
  assign ram_x_15_MPORT_addr = 1'h0;
  assign ram_x_15_MPORT_mask = 1'h1;
  assign ram_x_15_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_x_0 = ram_x_0_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_1 = ram_x_1_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_2 = ram_x_2_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_3 = ram_x_3_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_4 = ram_x_4_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_5 = ram_x_5_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_6 = ram_x_6_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_7 = ram_x_7_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_8 = ram_x_8_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_9 = ram_x_9_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_10 = ram_x_10_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_11 = ram_x_11_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_12 = ram_x_12_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_13 = ram_x_13_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_14 = ram_x_14_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_x_15 = ram_x_15_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_x_0_MPORT_en & ram_x_0_MPORT_mask) begin
      ram_x_0[ram_x_0_MPORT_addr] <= ram_x_0_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_1_MPORT_en & ram_x_1_MPORT_mask) begin
      ram_x_1[ram_x_1_MPORT_addr] <= ram_x_1_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_2_MPORT_en & ram_x_2_MPORT_mask) begin
      ram_x_2[ram_x_2_MPORT_addr] <= ram_x_2_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_3_MPORT_en & ram_x_3_MPORT_mask) begin
      ram_x_3[ram_x_3_MPORT_addr] <= ram_x_3_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_4_MPORT_en & ram_x_4_MPORT_mask) begin
      ram_x_4[ram_x_4_MPORT_addr] <= ram_x_4_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_5_MPORT_en & ram_x_5_MPORT_mask) begin
      ram_x_5[ram_x_5_MPORT_addr] <= ram_x_5_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_6_MPORT_en & ram_x_6_MPORT_mask) begin
      ram_x_6[ram_x_6_MPORT_addr] <= ram_x_6_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_7_MPORT_en & ram_x_7_MPORT_mask) begin
      ram_x_7[ram_x_7_MPORT_addr] <= ram_x_7_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_8_MPORT_en & ram_x_8_MPORT_mask) begin
      ram_x_8[ram_x_8_MPORT_addr] <= ram_x_8_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_9_MPORT_en & ram_x_9_MPORT_mask) begin
      ram_x_9[ram_x_9_MPORT_addr] <= ram_x_9_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_10_MPORT_en & ram_x_10_MPORT_mask) begin
      ram_x_10[ram_x_10_MPORT_addr] <= ram_x_10_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_11_MPORT_en & ram_x_11_MPORT_mask) begin
      ram_x_11[ram_x_11_MPORT_addr] <= ram_x_11_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_12_MPORT_en & ram_x_12_MPORT_mask) begin
      ram_x_12[ram_x_12_MPORT_addr] <= ram_x_12_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_13_MPORT_en & ram_x_13_MPORT_mask) begin
      ram_x_13[ram_x_13_MPORT_addr] <= ram_x_13_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_14_MPORT_en & ram_x_14_MPORT_mask) begin
      ram_x_14[ram_x_14_MPORT_addr] <= ram_x_14_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_x_15_MPORT_en & ram_x_15_MPORT_mask) begin
      ram_x_15[ram_x_15_MPORT_addr] <= ram_x_15_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Decoupled.scala 279:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 280:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 262:27]
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_0[initvar] = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_1[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_2[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_3[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_4[initvar] = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_5[initvar] = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_6[initvar] = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_7[initvar] = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_8[initvar] = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_9[initvar] = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_10[initvar] = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_11[initvar] = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_12[initvar] = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_13[initvar] = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_14[initvar] = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_x_15[initvar] = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_16[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  maybe_full = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    maybe_full = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineHsk_1(
  input   clock,
  input   reset,
  input   io_validPre,
  output  io_readyPre,
  input   io_lastPre,
  output  io_validNxt,
  input   io_readyNxt,
  output  io_regen_0,
  output  io_lastNxt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  valid_1_r; // @[Reg.scala 28:20]
  wire  ready_0 = io_readyNxt | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  reg  last_1_r; // @[Reg.scala 28:20]
  assign io_readyPre = io_readyNxt | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  assign io_validNxt = valid_1_r; // @[pipelinehsk.scala 17:21 22:20]
  assign io_regen_0 = io_validPre & ready_0; // @[pipelinehsk.scala 25:33]
  assign io_lastNxt = last_1_r; // @[pipelinehsk.scala 19:20 23:19]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_0) begin // @[Reg.scala 28:20]
      valid_1_r <= io_validPre;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_0) begin // @[Reg.scala 28:20]
      last_1_r <= io_lastPre;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_1_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  last_1_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid_1_r = 1'h0;
  end
  if (reset) begin
    last_1_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Adder2to1(
  input        clock,
  input        reset,
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_x_0,
  input  [7:0] io_input_bits_x_1,
  input  [7:0] io_input_bits_x_2,
  input  [7:0] io_input_bits_x_3,
  input  [7:0] io_input_bits_x_4,
  input  [7:0] io_input_bits_x_5,
  input  [7:0] io_input_bits_x_6,
  input  [7:0] io_input_bits_x_7,
  input  [7:0] io_input_bits_x_8,
  input  [7:0] io_input_bits_x_9,
  input  [7:0] io_input_bits_x_10,
  input  [7:0] io_input_bits_x_11,
  input  [7:0] io_input_bits_x_12,
  input  [7:0] io_input_bits_x_13,
  input  [7:0] io_input_bits_x_14,
  input  [7:0] io_input_bits_x_15,
  input  [7:0] io_input_bits_x_16,
  input  [7:0] io_input_bits_x_17,
  input  [7:0] io_input_bits_x_18,
  input  [7:0] io_input_bits_x_19,
  input  [7:0] io_input_bits_x_20,
  input  [7:0] io_input_bits_x_21,
  input  [7:0] io_input_bits_x_22,
  input  [7:0] io_input_bits_x_23,
  input  [7:0] io_input_bits_x_24,
  input  [7:0] io_input_bits_x_25,
  input  [7:0] io_input_bits_x_26,
  input  [7:0] io_input_bits_x_27,
  input  [7:0] io_input_bits_x_28,
  input  [7:0] io_input_bits_x_29,
  input  [7:0] io_input_bits_x_30,
  input  [7:0] io_input_bits_x_31,
  input        io_input_bits_last,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_x_0,
  output [7:0] io_output_bits_x_1,
  output [7:0] io_output_bits_x_2,
  output [7:0] io_output_bits_x_3,
  output [7:0] io_output_bits_x_4,
  output [7:0] io_output_bits_x_5,
  output [7:0] io_output_bits_x_6,
  output [7:0] io_output_bits_x_7,
  output [7:0] io_output_bits_x_8,
  output [7:0] io_output_bits_x_9,
  output [7:0] io_output_bits_x_10,
  output [7:0] io_output_bits_x_11,
  output [7:0] io_output_bits_x_12,
  output [7:0] io_output_bits_x_13,
  output [7:0] io_output_bits_x_14,
  output [7:0] io_output_bits_x_15,
  output       io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  hsk_clock; // @[adder2to1.scala 26:25]
  wire  hsk_reset; // @[adder2to1.scala 26:25]
  wire  hsk_io_validPre; // @[adder2to1.scala 26:25]
  wire  hsk_io_readyPre; // @[adder2to1.scala 26:25]
  wire  hsk_io_lastPre; // @[adder2to1.scala 26:25]
  wire  hsk_io_validNxt; // @[adder2to1.scala 26:25]
  wire  hsk_io_readyNxt; // @[adder2to1.scala 26:25]
  wire  hsk_io_regen_0; // @[adder2to1.scala 26:25]
  wire  hsk_io_lastNxt; // @[adder2to1.scala 26:25]
  wire [7:0] sum_0 = $signed(io_input_bits_x_0) + $signed(io_input_bits_x_16); // @[adder2to1.scala 23:69]
  wire [7:0] sum_1 = $signed(io_input_bits_x_1) + $signed(io_input_bits_x_17); // @[adder2to1.scala 23:69]
  wire [7:0] sum_2 = $signed(io_input_bits_x_2) + $signed(io_input_bits_x_18); // @[adder2to1.scala 23:69]
  wire [7:0] sum_3 = $signed(io_input_bits_x_3) + $signed(io_input_bits_x_19); // @[adder2to1.scala 23:69]
  wire [7:0] sum_4 = $signed(io_input_bits_x_4) + $signed(io_input_bits_x_20); // @[adder2to1.scala 23:69]
  wire [7:0] sum_5 = $signed(io_input_bits_x_5) + $signed(io_input_bits_x_21); // @[adder2to1.scala 23:69]
  wire [7:0] sum_6 = $signed(io_input_bits_x_6) + $signed(io_input_bits_x_22); // @[adder2to1.scala 23:69]
  wire [7:0] sum_7 = $signed(io_input_bits_x_7) + $signed(io_input_bits_x_23); // @[adder2to1.scala 23:69]
  wire [7:0] sum_8 = $signed(io_input_bits_x_8) + $signed(io_input_bits_x_24); // @[adder2to1.scala 23:69]
  wire [7:0] sum_9 = $signed(io_input_bits_x_9) + $signed(io_input_bits_x_25); // @[adder2to1.scala 23:69]
  wire [7:0] sum_10 = $signed(io_input_bits_x_10) + $signed(io_input_bits_x_26); // @[adder2to1.scala 23:69]
  wire [7:0] sum_11 = $signed(io_input_bits_x_11) + $signed(io_input_bits_x_27); // @[adder2to1.scala 23:69]
  wire [7:0] sum_12 = $signed(io_input_bits_x_12) + $signed(io_input_bits_x_28); // @[adder2to1.scala 23:69]
  wire [7:0] sum_13 = $signed(io_input_bits_x_13) + $signed(io_input_bits_x_29); // @[adder2to1.scala 23:69]
  wire [7:0] sum_14 = $signed(io_input_bits_x_14) + $signed(io_input_bits_x_30); // @[adder2to1.scala 23:69]
  wire [7:0] sum_15 = $signed(io_input_bits_x_15) + $signed(io_input_bits_x_31); // @[adder2to1.scala 23:69]
  reg [7:0] r_0; // @[Reg.scala 16:16]
  reg [7:0] r_1; // @[Reg.scala 16:16]
  reg [7:0] r_2; // @[Reg.scala 16:16]
  reg [7:0] r_3; // @[Reg.scala 16:16]
  reg [7:0] r_4; // @[Reg.scala 16:16]
  reg [7:0] r_5; // @[Reg.scala 16:16]
  reg [7:0] r_6; // @[Reg.scala 16:16]
  reg [7:0] r_7; // @[Reg.scala 16:16]
  reg [7:0] r_8; // @[Reg.scala 16:16]
  reg [7:0] r_9; // @[Reg.scala 16:16]
  reg [7:0] r_10; // @[Reg.scala 16:16]
  reg [7:0] r_11; // @[Reg.scala 16:16]
  reg [7:0] r_12; // @[Reg.scala 16:16]
  reg [7:0] r_13; // @[Reg.scala 16:16]
  reg [7:0] r_14; // @[Reg.scala 16:16]
  reg [7:0] r_15; // @[Reg.scala 16:16]
  PipelineHsk_1 hsk ( // @[adder2to1.scala 26:25]
    .clock(hsk_clock),
    .reset(hsk_reset),
    .io_validPre(hsk_io_validPre),
    .io_readyPre(hsk_io_readyPre),
    .io_lastPre(hsk_io_lastPre),
    .io_validNxt(hsk_io_validNxt),
    .io_readyNxt(hsk_io_readyNxt),
    .io_regen_0(hsk_io_regen_0),
    .io_lastNxt(hsk_io_lastNxt)
  );
  assign io_input_ready = hsk_io_readyPre; // @[adder2to1.scala 28:24]
  assign io_output_valid = hsk_io_validNxt; // @[adder2to1.scala 29:25]
  assign io_output_bits_x_0 = r_0; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_1 = r_1; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_2 = r_2; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_3 = r_3; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_4 = r_4; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_5 = r_5; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_6 = r_6; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_7 = r_7; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_8 = r_8; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_9 = r_9; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_10 = r_10; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_11 = r_11; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_12 = r_12; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_13 = r_13; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_14 = r_14; // @[adder2to1.scala 33:26]
  assign io_output_bits_x_15 = r_15; // @[adder2to1.scala 33:26]
  assign io_output_bits_last = hsk_io_lastNxt; // @[adder2to1.scala 32:29]
  assign hsk_clock = clock;
  assign hsk_reset = reset;
  assign hsk_io_validPre = io_input_valid; // @[adder2to1.scala 27:25]
  assign hsk_io_lastPre = io_input_bits_last; // @[adder2to1.scala 31:24]
  assign hsk_io_readyNxt = io_output_ready; // @[adder2to1.scala 30:25]
  always @(posedge clock) begin
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_0 <= sum_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_1 <= sum_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_2 <= sum_2; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_3 <= sum_3; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_4 <= sum_4; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_5 <= sum_5; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_6 <= sum_6; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_7 <= sum_7; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_8 <= sum_8; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_9 <= sum_9; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_10 <= sum_10; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_11 <= sum_11; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_12 <= sum_12; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_13 <= sum_13; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_14 <= sum_14; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_15 <= sum_15; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  r_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  r_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  r_15 = _RAND_15[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineHsk_2(
  input   clock,
  input   reset,
  input   io_validPre,
  output  io_readyPre,
  input   io_lastPre,
  output  io_validNxt,
  input   io_readyNxt,
  output  io_regen_0,
  output  io_regen_1,
  output  io_regen_2,
  output  io_regen_3,
  output  io_lastNxt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  valid_1_r; // @[Reg.scala 28:20]
  reg  valid_4_r; // @[Reg.scala 28:20]
  wire  ready_3 = io_readyNxt | ~valid_4_r; // @[pipelinehsk.scala 24:32]
  reg  valid_3_r; // @[Reg.scala 28:20]
  wire  ready_2 = ready_3 | ~valid_3_r; // @[pipelinehsk.scala 24:32]
  reg  valid_2_r; // @[Reg.scala 28:20]
  wire  ready_1 = ready_2 | ~valid_2_r; // @[pipelinehsk.scala 24:32]
  wire  ready_0 = ready_1 | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  reg  last_1_r; // @[Reg.scala 28:20]
  reg  last_2_r; // @[Reg.scala 28:20]
  reg  last_3_r; // @[Reg.scala 28:20]
  reg  last_4_r; // @[Reg.scala 28:20]
  assign io_readyPre = ready_1 | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  assign io_validNxt = valid_4_r; // @[pipelinehsk.scala 17:21 22:20]
  assign io_regen_0 = io_validPre & ready_0; // @[pipelinehsk.scala 25:33]
  assign io_regen_1 = valid_1_r & ready_1; // @[pipelinehsk.scala 25:33]
  assign io_regen_2 = valid_2_r & ready_2; // @[pipelinehsk.scala 25:33]
  assign io_regen_3 = valid_3_r & ready_3; // @[pipelinehsk.scala 25:33]
  assign io_lastNxt = last_4_r; // @[pipelinehsk.scala 19:20 23:19]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_0) begin // @[Reg.scala 28:20]
      valid_1_r <= io_validPre;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_4_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_3) begin // @[Reg.scala 28:20]
      valid_4_r <= valid_3_r;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_3_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_2) begin // @[Reg.scala 28:20]
      valid_3_r <= valid_2_r;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_2_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_1) begin // @[Reg.scala 28:20]
      valid_2_r <= valid_1_r;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_0) begin // @[Reg.scala 28:20]
      last_1_r <= io_lastPre;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_2_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_1) begin // @[Reg.scala 28:20]
      last_2_r <= last_1_r;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_3_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_2) begin // @[Reg.scala 28:20]
      last_3_r <= last_2_r;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_4_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_3) begin // @[Reg.scala 28:20]
      last_4_r <= last_3_r;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_1_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_4_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_3_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_2_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  last_1_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  last_2_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  last_3_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  last_4_r = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid_1_r = 1'h0;
  end
  if (reset) begin
    valid_4_r = 1'h0;
  end
  if (reset) begin
    valid_3_r = 1'h0;
  end
  if (reset) begin
    valid_2_r = 1'h0;
  end
  if (reset) begin
    last_1_r = 1'h0;
  end
  if (reset) begin
    last_2_r = 1'h0;
  end
  if (reset) begin
    last_3_r = 1'h0;
  end
  if (reset) begin
    last_4_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AdderTree(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [11:0] io_input_bits_x_0,
  input  [11:0] io_input_bits_x_1,
  input  [11:0] io_input_bits_x_2,
  input  [11:0] io_input_bits_x_3,
  input  [11:0] io_input_bits_x_4,
  input  [11:0] io_input_bits_x_5,
  input  [11:0] io_input_bits_x_6,
  input  [11:0] io_input_bits_x_7,
  input  [11:0] io_input_bits_x_8,
  input  [11:0] io_input_bits_x_9,
  input  [11:0] io_input_bits_x_10,
  input  [11:0] io_input_bits_x_11,
  input  [11:0] io_input_bits_x_12,
  input  [11:0] io_input_bits_x_13,
  input  [11:0] io_input_bits_x_14,
  input  [11:0] io_input_bits_x_15,
  input         io_input_bits_last,
  output        io_output_valid,
  output [11:0] io_output_bits_x_0,
  output        io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  hsk_clock; // @[addertree.scala 32:21]
  wire  hsk_reset; // @[addertree.scala 32:21]
  wire  hsk_io_validPre; // @[addertree.scala 32:21]
  wire  hsk_io_readyPre; // @[addertree.scala 32:21]
  wire  hsk_io_lastPre; // @[addertree.scala 32:21]
  wire  hsk_io_validNxt; // @[addertree.scala 32:21]
  wire  hsk_io_readyNxt; // @[addertree.scala 32:21]
  wire  hsk_io_regen_0; // @[addertree.scala 32:21]
  wire  hsk_io_regen_1; // @[addertree.scala 32:21]
  wire  hsk_io_regen_2; // @[addertree.scala 32:21]
  wire  hsk_io_regen_3; // @[addertree.scala 32:21]
  wire  hsk_io_lastNxt; // @[addertree.scala 32:21]
  reg [11:0] r; // @[Reg.scala 16:16]
  wire [11:0] _s_T_2 = io_input_bits_x_0 ^ io_input_bits_x_4; // @[addertree.scala 72:46]
  wire [11:0] s = _s_T_2 ^ io_input_bits_x_8; // @[addertree.scala 72:80]
  wire [11:0] _c_T_2 = io_input_bits_x_0 & io_input_bits_x_4; // @[addertree.scala 73:46]
  wire [11:0] _c_T_5 = io_input_bits_x_0 & io_input_bits_x_8; // @[addertree.scala 73:108]
  wire [11:0] _c_T_6 = _c_T_2 | _c_T_5; // @[addertree.scala 73:80]
  wire [11:0] _c_T_9 = io_input_bits_x_4 & io_input_bits_x_8; // @[addertree.scala 73:178]
  wire [11:0] _c_T_10 = _c_T_6 | _c_T_9; // @[addertree.scala 73:144]
  wire [12:0] _c_T_11 = {_c_T_10, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c = _c_T_11[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_1_0_T = s ^ c; // @[addertree.scala 74:40]
  wire [11:0] sumIn_1_0 = _sumIn_1_0_T ^ io_input_bits_x_12; // @[addertree.scala 74:92]
  reg [11:0] r_1; // @[Reg.scala 16:16]
  wire [11:0] _s_T_7 = io_input_bits_x_1 ^ io_input_bits_x_5; // @[addertree.scala 72:46]
  wire [11:0] s_1 = _s_T_7 ^ io_input_bits_x_9; // @[addertree.scala 72:80]
  wire [11:0] _c_T_14 = io_input_bits_x_1 & io_input_bits_x_5; // @[addertree.scala 73:46]
  wire [11:0] _c_T_17 = io_input_bits_x_1 & io_input_bits_x_9; // @[addertree.scala 73:108]
  wire [11:0] _c_T_18 = _c_T_14 | _c_T_17; // @[addertree.scala 73:80]
  wire [11:0] _c_T_21 = io_input_bits_x_5 & io_input_bits_x_9; // @[addertree.scala 73:178]
  wire [11:0] _c_T_22 = _c_T_18 | _c_T_21; // @[addertree.scala 73:144]
  wire [12:0] _c_T_23 = {_c_T_22, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c_1 = _c_T_23[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_1_1_T = s_1 ^ c_1; // @[addertree.scala 74:40]
  wire [11:0] sumIn_1_1 = _sumIn_1_1_T ^ io_input_bits_x_13; // @[addertree.scala 74:92]
  reg [11:0] r_2; // @[Reg.scala 16:16]
  wire [11:0] _s_T_12 = io_input_bits_x_2 ^ io_input_bits_x_6; // @[addertree.scala 72:46]
  wire [11:0] s_2 = _s_T_12 ^ io_input_bits_x_10; // @[addertree.scala 72:80]
  wire [11:0] _c_T_26 = io_input_bits_x_2 & io_input_bits_x_6; // @[addertree.scala 73:46]
  wire [11:0] _c_T_29 = io_input_bits_x_2 & io_input_bits_x_10; // @[addertree.scala 73:108]
  wire [11:0] _c_T_30 = _c_T_26 | _c_T_29; // @[addertree.scala 73:80]
  wire [11:0] _c_T_33 = io_input_bits_x_6 & io_input_bits_x_10; // @[addertree.scala 73:178]
  wire [11:0] _c_T_34 = _c_T_30 | _c_T_33; // @[addertree.scala 73:144]
  wire [12:0] _c_T_35 = {_c_T_34, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c_2 = _c_T_35[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_1_2_T = s_2 ^ c_2; // @[addertree.scala 74:40]
  wire [11:0] sumIn_1_2 = _sumIn_1_2_T ^ io_input_bits_x_14; // @[addertree.scala 74:92]
  reg [11:0] r_3; // @[Reg.scala 16:16]
  wire [11:0] _s_T_17 = io_input_bits_x_3 ^ io_input_bits_x_7; // @[addertree.scala 72:46]
  wire [11:0] s_3 = _s_T_17 ^ io_input_bits_x_11; // @[addertree.scala 72:80]
  wire [11:0] _c_T_38 = io_input_bits_x_3 & io_input_bits_x_7; // @[addertree.scala 73:46]
  wire [11:0] _c_T_41 = io_input_bits_x_3 & io_input_bits_x_11; // @[addertree.scala 73:108]
  wire [11:0] _c_T_42 = _c_T_38 | _c_T_41; // @[addertree.scala 73:80]
  wire [11:0] _c_T_45 = io_input_bits_x_7 & io_input_bits_x_11; // @[addertree.scala 73:178]
  wire [11:0] _c_T_46 = _c_T_42 | _c_T_45; // @[addertree.scala 73:144]
  wire [12:0] _c_T_47 = {_c_T_46, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c_3 = _c_T_47[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_1_3_T = s_3 ^ c_3; // @[addertree.scala 74:40]
  wire [11:0] sumIn_1_3 = _sumIn_1_3_T ^ io_input_bits_x_15; // @[addertree.scala 74:92]
  reg [11:0] r_4; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_1_4_T = s & c; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_1_4_T_2 = s & io_input_bits_x_12; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_1_4_T_3 = _sumIn_1_4_T | _sumIn_1_4_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_1_4_T_5 = c & io_input_bits_x_12; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_1_4_T_7 = _sumIn_1_4_T_3 | _sumIn_1_4_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_1_4_T_8 = {$signed(_sumIn_1_4_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_1_4 = _sumIn_1_4_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_5; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_1_5_T = s_1 & c_1; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_1_5_T_2 = s_1 & io_input_bits_x_13; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_1_5_T_3 = _sumIn_1_5_T | _sumIn_1_5_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_1_5_T_5 = c_1 & io_input_bits_x_13; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_1_5_T_7 = _sumIn_1_5_T_3 | _sumIn_1_5_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_1_5_T_8 = {$signed(_sumIn_1_5_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_1_5 = _sumIn_1_5_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_6; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_1_6_T = s_2 & c_2; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_1_6_T_2 = s_2 & io_input_bits_x_14; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_1_6_T_3 = _sumIn_1_6_T | _sumIn_1_6_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_1_6_T_5 = c_2 & io_input_bits_x_14; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_1_6_T_7 = _sumIn_1_6_T_3 | _sumIn_1_6_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_1_6_T_8 = {$signed(_sumIn_1_6_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_1_6 = _sumIn_1_6_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_7; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_1_7_T = s_3 & c_3; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_1_7_T_2 = s_3 & io_input_bits_x_15; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_1_7_T_3 = _sumIn_1_7_T | _sumIn_1_7_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_1_7_T_5 = c_3 & io_input_bits_x_15; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_1_7_T_7 = _sumIn_1_7_T_3 | _sumIn_1_7_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_1_7_T_8 = {$signed(_sumIn_1_7_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_1_7 = _sumIn_1_7_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_16; // @[Reg.scala 16:16]
  wire [11:0] _s_T_22 = r ^ r_2; // @[addertree.scala 72:46]
  wire [11:0] s_4 = _s_T_22 ^ r_4; // @[addertree.scala 72:80]
  wire [11:0] _c_T_50 = r & r_2; // @[addertree.scala 73:46]
  wire [11:0] _c_T_53 = r & r_4; // @[addertree.scala 73:108]
  wire [11:0] _c_T_54 = _c_T_50 | _c_T_53; // @[addertree.scala 73:80]
  wire [11:0] _c_T_57 = r_2 & r_4; // @[addertree.scala 73:178]
  wire [11:0] _c_T_58 = _c_T_54 | _c_T_57; // @[addertree.scala 73:144]
  wire [12:0] _c_T_59 = {_c_T_58, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c_4 = _c_T_59[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_2_0_T = s_4 ^ c_4; // @[addertree.scala 74:40]
  wire [11:0] sumIn_2_0 = _sumIn_2_0_T ^ r_6; // @[addertree.scala 74:92]
  reg [11:0] r_17; // @[Reg.scala 16:16]
  wire [11:0] _s_T_27 = r_1 ^ r_3; // @[addertree.scala 72:46]
  wire [11:0] s_5 = _s_T_27 ^ r_5; // @[addertree.scala 72:80]
  wire [11:0] _c_T_62 = r_1 & r_3; // @[addertree.scala 73:46]
  wire [11:0] _c_T_65 = r_1 & r_5; // @[addertree.scala 73:108]
  wire [11:0] _c_T_66 = _c_T_62 | _c_T_65; // @[addertree.scala 73:80]
  wire [11:0] _c_T_69 = r_3 & r_5; // @[addertree.scala 73:178]
  wire [11:0] _c_T_70 = _c_T_66 | _c_T_69; // @[addertree.scala 73:144]
  wire [12:0] _c_T_71 = {_c_T_70, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c_5 = _c_T_71[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_2_1_T = s_5 ^ c_5; // @[addertree.scala 74:40]
  wire [11:0] sumIn_2_1 = _sumIn_2_1_T ^ r_7; // @[addertree.scala 74:92]
  reg [11:0] r_18; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_2_2_T = s_4 & c_4; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_2_2_T_2 = s_4 & r_6; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_2_2_T_3 = _sumIn_2_2_T | _sumIn_2_2_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_2_2_T_5 = c_4 & r_6; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_2_2_T_7 = _sumIn_2_2_T_3 | _sumIn_2_2_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_2_2_T_8 = {$signed(_sumIn_2_2_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_2_2 = _sumIn_2_2_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_19; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_2_3_T = s_5 & c_5; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_2_3_T_2 = s_5 & r_7; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_2_3_T_3 = _sumIn_2_3_T | _sumIn_2_3_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_2_3_T_5 = c_5 & r_7; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_2_3_T_7 = _sumIn_2_3_T_3 | _sumIn_2_3_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_2_3_T_8 = {$signed(_sumIn_2_3_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_2_3 = _sumIn_2_3_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_32; // @[Reg.scala 16:16]
  wire [11:0] _s_T_32 = r_16 ^ r_17; // @[addertree.scala 72:46]
  wire [11:0] s_6 = _s_T_32 ^ r_18; // @[addertree.scala 72:80]
  wire [11:0] _c_T_74 = r_16 & r_17; // @[addertree.scala 73:46]
  wire [11:0] _c_T_77 = r_16 & r_18; // @[addertree.scala 73:108]
  wire [11:0] _c_T_78 = _c_T_74 | _c_T_77; // @[addertree.scala 73:80]
  wire [11:0] _c_T_81 = r_17 & r_18; // @[addertree.scala 73:178]
  wire [11:0] _c_T_82 = _c_T_78 | _c_T_81; // @[addertree.scala 73:144]
  wire [12:0] _c_T_83 = {_c_T_82, 1'h0}; // @[addertree.scala 73:215]
  wire [11:0] c_6 = _c_T_83[11:0]; // @[addertree.scala 71:25 73:15]
  wire [11:0] _sumIn_3_0_T = s_6 ^ c_6; // @[addertree.scala 74:40]
  wire [11:0] sumIn_3_0 = _sumIn_3_0_T ^ r_19; // @[addertree.scala 74:92]
  reg [11:0] r_33; // @[Reg.scala 16:16]
  wire [11:0] _sumIn_3_1_T = s_6 & c_6; // @[addertree.scala 75:47]
  wire [11:0] _sumIn_3_1_T_2 = s_6 & r_19; // @[addertree.scala 75:53]
  wire [11:0] _sumIn_3_1_T_3 = _sumIn_3_1_T | _sumIn_3_1_T_2; // @[addertree.scala 75:50]
  wire [11:0] _sumIn_3_1_T_5 = c_6 & r_19; // @[addertree.scala 75:93]
  wire [11:0] _sumIn_3_1_T_7 = _sumIn_3_1_T_3 | _sumIn_3_1_T_5; // @[addertree.scala 75:143]
  wire [12:0] _sumIn_3_1_T_8 = {$signed(_sumIn_3_1_T_7), 1'h0}; // @[addertree.scala 75:154]
  wire [11:0] sumIn_3_1 = _sumIn_3_1_T_8[11:0]; // @[addertree.scala 41:21 75:41]
  reg [11:0] r_48; // @[Reg.scala 16:16]
  wire [11:0] sumIn_4_0 = $signed(r_32) + $signed(r_33); // @[addertree.scala 88:63]
  PipelineHsk_2 hsk ( // @[addertree.scala 32:21]
    .clock(hsk_clock),
    .reset(hsk_reset),
    .io_validPre(hsk_io_validPre),
    .io_readyPre(hsk_io_readyPre),
    .io_lastPre(hsk_io_lastPre),
    .io_validNxt(hsk_io_validNxt),
    .io_readyNxt(hsk_io_readyNxt),
    .io_regen_0(hsk_io_regen_0),
    .io_regen_1(hsk_io_regen_1),
    .io_regen_2(hsk_io_regen_2),
    .io_regen_3(hsk_io_regen_3),
    .io_lastNxt(hsk_io_lastNxt)
  );
  assign io_input_ready = hsk_io_readyPre; // @[addertree.scala 34:20]
  assign io_output_valid = hsk_io_validNxt; // @[addertree.scala 36:21]
  assign io_output_bits_x_0 = r_48; // @[addertree.scala 42:22 51:31]
  assign io_output_bits_last = hsk_io_lastNxt; // @[addertree.scala 38:25]
  assign hsk_clock = clock;
  assign hsk_reset = reset;
  assign hsk_io_validPre = io_input_valid; // @[addertree.scala 33:21]
  assign hsk_io_lastPre = io_input_bits_last; // @[addertree.scala 35:20]
  assign hsk_io_readyNxt = 1'h1; // @[addertree.scala 37:21]
  always @(posedge clock) begin
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r <= sumIn_1_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_1 <= sumIn_1_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_2 <= sumIn_1_2; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_3 <= sumIn_1_3; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_4 <= sumIn_1_4; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_5 <= sumIn_1_5; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_6 <= sumIn_1_6; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_7 <= sumIn_1_7; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      r_16 <= sumIn_2_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      r_17 <= sumIn_2_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      r_18 <= sumIn_2_2; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      r_19 <= sumIn_2_3; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_2) begin // @[Reg.scala 17:18]
      r_32 <= sumIn_3_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_2) begin // @[Reg.scala 17:18]
      r_33 <= sumIn_3_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_3) begin // @[Reg.scala 17:18]
      r_48 <= sumIn_4_0; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  r_6 = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  r_7 = _RAND_7[11:0];
  _RAND_8 = {1{`RANDOM}};
  r_16 = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  r_17 = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  r_18 = _RAND_10[11:0];
  _RAND_11 = {1{`RANDOM}};
  r_19 = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  r_32 = _RAND_12[11:0];
  _RAND_13 = {1{`RANDOM}};
  r_33 = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  r_48 = _RAND_14[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Accumulator2to1(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [11:0] io_input_bits_x_0,
  input         io_input_bits_last,
  output        io_output_valid,
  output [11:0] io_output_bits_x_0,
  output        io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _io_output_bits_last_T = io_input_valid & io_input_ready; // @[accumulator2to1.scala 17:77]
  reg  io_output_bits_last_r; // @[Reg.scala 28:20]
  reg [11:0] io_output_bits_x_0_r; // @[Reg.scala 28:20]
  wire [11:0] _sumNxt_T_2 = $signed(io_output_bits_x_0) + $signed(io_input_bits_x_0); // @[accumulator2to1.scala 19:79]
  assign io_input_ready = 1'h1; // @[accumulator2to1.scala 15:20]
  assign io_output_valid = io_output_bits_last; // @[accumulator2to1.scala 20:21]
  assign io_output_bits_x_0 = io_output_bits_x_0_r; // @[accumulator2to1.scala 18:25]
  assign io_output_bits_last = io_output_bits_last_r; // @[accumulator2to1.scala 17:25]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      io_output_bits_last_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (_io_output_bits_last_T) begin // @[Reg.scala 28:20]
      io_output_bits_last_r <= io_input_bits_last;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      io_output_bits_x_0_r <= 12'sh0; // @[accumulator2to1.scala 19:18]
    end else if (_io_output_bits_last_T) begin // @[Reg.scala 28:20]
      if (io_output_bits_last) begin
        io_output_bits_x_0_r <= io_input_bits_x_0;
      end else begin
        io_output_bits_x_0_r <= _sumNxt_T_2;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_output_bits_last_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_output_bits_x_0_r = _RAND_1[11:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    io_output_bits_last_r = 1'h0;
  end
  if (reset) begin
    io_output_bits_x_0_r = 12'sh0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Logarithm(
  input         clock,
  input         reset,
  input         io_input_valid,
  input  [11:0] io_input_bits_x_0,
  input         io_input_bits_last,
  input         io_output_ready,
  output        io_output_valid,
  output [7:0]  io_output_bits_x_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  hsk_clock; // @[logarithm.scala 19:21]
  wire  hsk_reset; // @[logarithm.scala 19:21]
  wire  hsk_io_validPre; // @[logarithm.scala 19:21]
  wire  hsk_io_readyPre; // @[logarithm.scala 19:21]
  wire  hsk_io_lastPre; // @[logarithm.scala 19:21]
  wire  hsk_io_validNxt; // @[logarithm.scala 19:21]
  wire  hsk_io_readyNxt; // @[logarithm.scala 19:21]
  wire  hsk_io_regen_0; // @[logarithm.scala 19:21]
  wire  hsk_io_regen_1; // @[logarithm.scala 19:21]
  wire  hsk_io_regen_2; // @[logarithm.scala 19:21]
  wire  hsk_io_regen_3; // @[logarithm.scala 19:21]
  wire  hsk_io_lastNxt; // @[logarithm.scala 19:21]
  wire  lod_0_12 = io_input_bits_x_0[11]; // @[logarithm.scala 30:43]
  wire  lod_0_0 = $signed(io_input_bits_x_0) == 12'sh0; // @[logarithm.scala 31:40]
  wire  lod_0_1 = ~(io_input_bits_x_0[1] | io_input_bits_x_0[2] | io_input_bits_x_0[3] | io_input_bits_x_0[4] |
    io_input_bits_x_0[5] | io_input_bits_x_0[6] | io_input_bits_x_0[7] | io_input_bits_x_0[8] | io_input_bits_x_0[9] |
    io_input_bits_x_0[10] | io_input_bits_x_0[11]) & io_input_bits_x_0[0]; // @[logarithm.scala 33:83]
  wire  lod_0_2 = ~(io_input_bits_x_0[2] | io_input_bits_x_0[3] | io_input_bits_x_0[4] | io_input_bits_x_0[5] |
    io_input_bits_x_0[6] | io_input_bits_x_0[7] | io_input_bits_x_0[8] | io_input_bits_x_0[9] | io_input_bits_x_0[10] |
    io_input_bits_x_0[11]) & io_input_bits_x_0[1]; // @[logarithm.scala 33:83]
  wire  lod_0_3 = ~(io_input_bits_x_0[3] | io_input_bits_x_0[4] | io_input_bits_x_0[5] | io_input_bits_x_0[6] |
    io_input_bits_x_0[7] | io_input_bits_x_0[8] | io_input_bits_x_0[9] | io_input_bits_x_0[10] | io_input_bits_x_0[11])
     & io_input_bits_x_0[2]; // @[logarithm.scala 33:83]
  wire  lod_0_4 = ~(io_input_bits_x_0[4] | io_input_bits_x_0[5] | io_input_bits_x_0[6] | io_input_bits_x_0[7] |
    io_input_bits_x_0[8] | io_input_bits_x_0[9] | io_input_bits_x_0[10] | io_input_bits_x_0[11]) & io_input_bits_x_0[3]; // @[logarithm.scala 33:83]
  wire  lod_0_5 = ~(io_input_bits_x_0[5] | io_input_bits_x_0[6] | io_input_bits_x_0[7] | io_input_bits_x_0[8] |
    io_input_bits_x_0[9] | io_input_bits_x_0[10] | io_input_bits_x_0[11]) & io_input_bits_x_0[4]; // @[logarithm.scala 33:83]
  wire  lod_0_6 = ~(io_input_bits_x_0[6] | io_input_bits_x_0[7] | io_input_bits_x_0[8] | io_input_bits_x_0[9] |
    io_input_bits_x_0[10] | io_input_bits_x_0[11]) & io_input_bits_x_0[5]; // @[logarithm.scala 33:83]
  wire  lod_0_7 = ~(io_input_bits_x_0[7] | io_input_bits_x_0[8] | io_input_bits_x_0[9] | io_input_bits_x_0[10] |
    io_input_bits_x_0[11]) & io_input_bits_x_0[6]; // @[logarithm.scala 33:83]
  wire  lod_0_8 = ~(io_input_bits_x_0[8] | io_input_bits_x_0[9] | io_input_bits_x_0[10] | io_input_bits_x_0[11]) &
    io_input_bits_x_0[7]; // @[logarithm.scala 33:83]
  wire  lod_0_9 = ~(io_input_bits_x_0[9] | io_input_bits_x_0[10] | io_input_bits_x_0[11]) & io_input_bits_x_0[8]; // @[logarithm.scala 33:83]
  wire  lod_0_10 = ~(io_input_bits_x_0[10] | io_input_bits_x_0[11]) & io_input_bits_x_0[9]; // @[logarithm.scala 33:83]
  wire  lod_0_11 = ~lod_0_12 & io_input_bits_x_0[10]; // @[logarithm.scala 33:83]
  reg  data1Lod_0_0; // @[Reg.scala 16:16]
  reg  data1Lod_0_1; // @[Reg.scala 16:16]
  reg  data1Lod_0_2; // @[Reg.scala 16:16]
  reg  data1Lod_0_3; // @[Reg.scala 16:16]
  reg  data1Lod_0_4; // @[Reg.scala 16:16]
  reg  data1Lod_0_5; // @[Reg.scala 16:16]
  reg  data1Lod_0_6; // @[Reg.scala 16:16]
  reg  data1Lod_0_7; // @[Reg.scala 16:16]
  reg  data1Lod_0_8; // @[Reg.scala 16:16]
  reg  data1Lod_0_9; // @[Reg.scala 16:16]
  reg  data1Lod_0_10; // @[Reg.scala 16:16]
  reg  data1Lod_0_11; // @[Reg.scala 16:16]
  reg  data1Lod_0_12; // @[Reg.scala 16:16]
  reg [11:0] data1In_0; // @[Reg.scala 16:16]
  wire [23:0] _data2InMux_0_T = {$signed(data1In_0), 12'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_2 = data1Lod_0_0 ? _data2InMux_0_T[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [22:0] _data2InMux_0_T_3 = {$signed(data1In_0), 11'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_5 = data1Lod_0_1 ? _data2InMux_0_T_3[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [21:0] _data2InMux_0_T_6 = {$signed(data1In_0), 10'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_8 = data1Lod_0_2 ? _data2InMux_0_T_6[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [20:0] _data2InMux_0_T_9 = {$signed(data1In_0), 9'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_11 = data1Lod_0_3 ? _data2InMux_0_T_9[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [19:0] _data2InMux_0_T_12 = {$signed(data1In_0), 8'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_14 = data1Lod_0_4 ? _data2InMux_0_T_12[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [18:0] _data2InMux_0_T_15 = {$signed(data1In_0), 7'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_17 = data1Lod_0_5 ? _data2InMux_0_T_15[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [17:0] _data2InMux_0_T_18 = {$signed(data1In_0), 6'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_20 = data1Lod_0_6 ? _data2InMux_0_T_18[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [16:0] _data2InMux_0_T_21 = {$signed(data1In_0), 5'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_23 = data1Lod_0_7 ? _data2InMux_0_T_21[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [15:0] _data2InMux_0_T_24 = {$signed(data1In_0), 4'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_26 = data1Lod_0_8 ? _data2InMux_0_T_24[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [14:0] _data2InMux_0_T_27 = {$signed(data1In_0), 3'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_29 = data1Lod_0_9 ? _data2InMux_0_T_27[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [13:0] _data2InMux_0_T_30 = {$signed(data1In_0), 2'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_32 = data1Lod_0_10 ? _data2InMux_0_T_30[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [12:0] _data2InMux_0_T_33 = {$signed(data1In_0), 1'h0}; // @[logarithm.scala 43:52]
  wire [11:0] _data2InMux_0_T_35 = data1Lod_0_11 ? _data2InMux_0_T_33[11:0] : 12'h0; // @[logarithm.scala 43:37]
  wire [11:0] _data2InMux_0_T_38 = data1Lod_0_12 ? data1In_0 : 12'h0; // @[logarithm.scala 43:37]
  wire [11:0] _data2InMux_0_T_40 = _data2InMux_0_T_2 | _data2InMux_0_T_5; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_41 = _data2InMux_0_T_40 | _data2InMux_0_T_8; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_42 = _data2InMux_0_T_41 | _data2InMux_0_T_11; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_43 = _data2InMux_0_T_42 | _data2InMux_0_T_14; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_44 = _data2InMux_0_T_43 | _data2InMux_0_T_17; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_45 = _data2InMux_0_T_44 | _data2InMux_0_T_20; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_46 = _data2InMux_0_T_45 | _data2InMux_0_T_23; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_47 = _data2InMux_0_T_46 | _data2InMux_0_T_26; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_48 = _data2InMux_0_T_47 | _data2InMux_0_T_29; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_49 = _data2InMux_0_T_48 | _data2InMux_0_T_32; // @[logarithm.scala 44:33]
  wire [11:0] _data2InMux_0_T_50 = _data2InMux_0_T_49 | _data2InMux_0_T_35; // @[logarithm.scala 44:33]
  wire [11:0] data2InMux_0 = _data2InMux_0_T_50 | _data2InMux_0_T_38; // @[logarithm.scala 44:50]
  wire [4:0] _T_1 = data1Lod_0_1 ? $signed(-5'sh6) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_2 = data1Lod_0_2 ? $signed(-5'sh5) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_3 = data1Lod_0_3 ? $signed(-5'sh4) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_4 = data1Lod_0_4 ? $signed(-5'sh3) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_5 = data1Lod_0_5 ? $signed(-5'sh2) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_6 = data1Lod_0_6 ? $signed(-5'sh1) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_8 = data1Lod_0_8 ? $signed(5'sh1) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_9 = data1Lod_0_9 ? $signed(5'sh2) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_10 = data1Lod_0_10 ? $signed(5'sh3) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_11 = data1Lod_0_11 ? $signed(5'sh4) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_12 = data1Lod_0_12 ? $signed(5'sh5) : $signed(5'sh0); // @[logarithm.scala 46:33]
  wire [4:0] _T_14 = data1Lod_0_0 ? $signed(-5'sh7) : $signed(5'sh0); // @[logarithm.scala 47:36]
  wire [4:0] _T_16 = $signed(_T_14) | $signed(_T_1); // @[logarithm.scala 47:36]
  wire [4:0] _T_18 = $signed(_T_16) | $signed(_T_2); // @[logarithm.scala 47:36]
  wire [4:0] _T_20 = $signed(_T_18) | $signed(_T_3); // @[logarithm.scala 47:36]
  wire [4:0] _T_22 = $signed(_T_20) | $signed(_T_4); // @[logarithm.scala 47:36]
  wire [4:0] _T_24 = $signed(_T_22) | $signed(_T_5); // @[logarithm.scala 47:36]
  wire [4:0] _T_28 = $signed(_T_24) | $signed(_T_6); // @[logarithm.scala 47:36]
  wire [4:0] _T_30 = $signed(_T_28) | $signed(_T_8); // @[logarithm.scala 47:36]
  wire [4:0] _T_32 = $signed(_T_30) | $signed(_T_9); // @[logarithm.scala 47:36]
  wire [4:0] _T_34 = $signed(_T_32) | $signed(_T_10); // @[logarithm.scala 47:36]
  wire [4:0] _T_36 = $signed(_T_34) | $signed(_T_11); // @[logarithm.scala 47:36]
  wire [4:0] data2CountMux_0 = $signed(_T_36) | $signed(_T_12); // @[logarithm.scala 47:36]
  reg [11:0] data2In_0; // @[Reg.scala 16:16]
  reg [4:0] data2Count_0; // @[Reg.scala 16:16]
  reg [4:0] data3In1_0; // @[Reg.scala 16:16]
  wire [4:0] _GEN_82 = 11'h42 == data2In_0[10:0] ? $signed(5'sh1) : $signed(5'sh0); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_83 = 11'h43 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_82); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_84 = 11'h44 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_83); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_85 = 11'h45 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_84); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_86 = 11'h46 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_85); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_87 = 11'h47 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_86); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_88 = 11'h48 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_87); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_89 = 11'h49 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_88); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_90 = 11'h4a == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_89); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_91 = 11'h4b == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_90); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_92 = 11'h4c == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_91); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_93 = 11'h4d == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_92); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_94 = 11'h4e == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_93); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_95 = 11'h4f == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_94); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_96 = 11'h50 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_95); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_97 = 11'h51 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_96); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_98 = 11'h52 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_97); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_99 = 11'h53 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_98); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_100 = 11'h54 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_99); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_101 = 11'h55 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_100); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_102 = 11'h56 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_101); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_103 = 11'h57 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_102); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_104 = 11'h58 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_103); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_105 = 11'h59 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_104); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_106 = 11'h5a == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_105); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_107 = 11'h5b == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_106); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_108 = 11'h5c == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_107); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_109 = 11'h5d == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_108); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_110 = 11'h5e == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_109); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_111 = 11'h5f == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_110); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_112 = 11'h60 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_111); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_113 = 11'h61 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_112); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_114 = 11'h62 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_113); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_115 = 11'h63 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_114); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_116 = 11'h64 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_115); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_117 = 11'h65 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_116); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_118 = 11'h66 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_117); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_119 = 11'h67 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_118); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_120 = 11'h68 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_119); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_121 = 11'h69 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_120); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_122 = 11'h6a == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_121); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_123 = 11'h6b == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_122); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_124 = 11'h6c == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_123); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_125 = 11'h6d == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_124); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_126 = 11'h6e == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_125); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_127 = 11'h6f == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_126); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_128 = 11'h70 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_127); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_129 = 11'h71 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_128); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_130 = 11'h72 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_129); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_131 = 11'h73 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_130); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_132 = 11'h74 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_131); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_133 = 11'h75 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_132); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_134 = 11'h76 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_133); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_135 = 11'h77 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_134); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_136 = 11'h78 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_135); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_137 = 11'h79 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_136); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_138 = 11'h7a == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_137); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_139 = 11'h7b == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_138); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_140 = 11'h7c == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_139); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_141 = 11'h7d == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_140); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_142 = 11'h7e == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_141); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_143 = 11'h7f == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_142); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_144 = 11'h80 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_143); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_145 = 11'h81 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_144); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_146 = 11'h82 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_145); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_147 = 11'h83 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_146); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_148 = 11'h84 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_147); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_149 = 11'h85 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_148); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_150 = 11'h86 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_149); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_151 = 11'h87 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_150); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_152 = 11'h88 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_151); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_153 = 11'h89 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_152); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_154 = 11'h8a == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_153); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_155 = 11'h8b == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_154); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_156 = 11'h8c == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_155); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_157 = 11'h8d == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_156); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_158 = 11'h8e == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_157); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_159 = 11'h8f == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_158); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_160 = 11'h90 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_159); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_161 = 11'h91 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_160); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_162 = 11'h92 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_161); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_163 = 11'h93 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_162); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_164 = 11'h94 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_163); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_165 = 11'h95 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_164); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_166 = 11'h96 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_165); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_167 = 11'h97 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_166); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_168 = 11'h98 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_167); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_169 = 11'h99 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_168); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_170 = 11'h9a == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_169); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_171 = 11'h9b == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_170); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_172 = 11'h9c == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_171); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_173 = 11'h9d == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_172); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_174 = 11'h9e == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_173); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_175 = 11'h9f == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_174); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_176 = 11'ha0 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_175); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_177 = 11'ha1 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_176); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_178 = 11'ha2 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_177); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_179 = 11'ha3 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_178); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_180 = 11'ha4 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_179); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_181 = 11'ha5 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_180); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_182 = 11'ha6 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_181); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_183 = 11'ha7 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_182); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_184 = 11'ha8 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_183); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_185 = 11'ha9 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_184); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_186 = 11'haa == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_185); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_187 = 11'hab == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_186); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_188 = 11'hac == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_187); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_189 = 11'had == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_188); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_190 = 11'hae == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_189); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_191 = 11'haf == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_190); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_192 = 11'hb0 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_191); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_193 = 11'hb1 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_192); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_194 = 11'hb2 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_193); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_195 = 11'hb3 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_194); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_196 = 11'hb4 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_195); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_197 = 11'hb5 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_196); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_198 = 11'hb6 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_197); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_199 = 11'hb7 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_198); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_200 = 11'hb8 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_199); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_201 = 11'hb9 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_200); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_202 = 11'hba == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_201); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_203 = 11'hbb == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_202); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_204 = 11'hbc == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_203); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_205 = 11'hbd == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_204); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_206 = 11'hbe == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_205); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_207 = 11'hbf == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_206); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_208 = 11'hc0 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_207); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_209 = 11'hc1 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_208); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_210 = 11'hc2 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_209); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_211 = 11'hc3 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_210); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_212 = 11'hc4 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_211); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_213 = 11'hc5 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_212); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_214 = 11'hc6 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_213); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_215 = 11'hc7 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_214); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_216 = 11'hc8 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_215); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_217 = 11'hc9 == data2In_0[10:0] ? $signed(5'sh1) : $signed(_GEN_216); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_218 = 11'hca == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_217); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_219 = 11'hcb == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_218); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_220 = 11'hcc == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_219); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_221 = 11'hcd == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_220); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_222 = 11'hce == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_221); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_223 = 11'hcf == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_222); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_224 = 11'hd0 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_223); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_225 = 11'hd1 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_224); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_226 = 11'hd2 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_225); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_227 = 11'hd3 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_226); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_228 = 11'hd4 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_227); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_229 = 11'hd5 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_228); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_230 = 11'hd6 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_229); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_231 = 11'hd7 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_230); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_232 = 11'hd8 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_231); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_233 = 11'hd9 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_232); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_234 = 11'hda == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_233); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_235 = 11'hdb == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_234); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_236 = 11'hdc == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_235); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_237 = 11'hdd == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_236); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_238 = 11'hde == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_237); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_239 = 11'hdf == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_238); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_240 = 11'he0 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_239); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_241 = 11'he1 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_240); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_242 = 11'he2 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_241); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_243 = 11'he3 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_242); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_244 = 11'he4 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_243); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_245 = 11'he5 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_244); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_246 = 11'he6 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_245); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_247 = 11'he7 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_246); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_248 = 11'he8 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_247); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_249 = 11'he9 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_248); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_250 = 11'hea == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_249); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_251 = 11'heb == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_250); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_252 = 11'hec == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_251); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_253 = 11'hed == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_252); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_254 = 11'hee == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_253); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_255 = 11'hef == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_254); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_256 = 11'hf0 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_255); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_257 = 11'hf1 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_256); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_258 = 11'hf2 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_257); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_259 = 11'hf3 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_258); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_260 = 11'hf4 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_259); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_261 = 11'hf5 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_260); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_262 = 11'hf6 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_261); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_263 = 11'hf7 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_262); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_264 = 11'hf8 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_263); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_265 = 11'hf9 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_264); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_266 = 11'hfa == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_265); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_267 = 11'hfb == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_266); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_268 = 11'hfc == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_267); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_269 = 11'hfd == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_268); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_270 = 11'hfe == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_269); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_271 = 11'hff == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_270); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_272 = 11'h100 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_271); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_273 = 11'h101 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_272); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_274 = 11'h102 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_273); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_275 = 11'h103 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_274); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_276 = 11'h104 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_275); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_277 = 11'h105 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_276); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_278 = 11'h106 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_277); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_279 = 11'h107 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_278); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_280 = 11'h108 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_279); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_281 = 11'h109 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_280); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_282 = 11'h10a == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_281); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_283 = 11'h10b == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_282); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_284 = 11'h10c == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_283); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_285 = 11'h10d == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_284); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_286 = 11'h10e == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_285); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_287 = 11'h10f == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_286); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_288 = 11'h110 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_287); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_289 = 11'h111 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_288); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_290 = 11'h112 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_289); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_291 = 11'h113 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_290); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_292 = 11'h114 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_291); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_293 = 11'h115 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_292); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_294 = 11'h116 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_293); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_295 = 11'h117 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_294); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_296 = 11'h118 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_295); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_297 = 11'h119 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_296); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_298 = 11'h11a == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_297); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_299 = 11'h11b == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_298); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_300 = 11'h11c == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_299); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_301 = 11'h11d == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_300); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_302 = 11'h11e == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_301); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_303 = 11'h11f == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_302); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_304 = 11'h120 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_303); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_305 = 11'h121 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_304); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_306 = 11'h122 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_305); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_307 = 11'h123 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_306); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_308 = 11'h124 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_307); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_309 = 11'h125 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_308); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_310 = 11'h126 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_309); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_311 = 11'h127 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_310); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_312 = 11'h128 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_311); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_313 = 11'h129 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_312); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_314 = 11'h12a == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_313); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_315 = 11'h12b == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_314); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_316 = 11'h12c == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_315); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_317 = 11'h12d == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_316); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_318 = 11'h12e == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_317); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_319 = 11'h12f == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_318); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_320 = 11'h130 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_319); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_321 = 11'h131 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_320); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_322 = 11'h132 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_321); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_323 = 11'h133 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_322); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_324 = 11'h134 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_323); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_325 = 11'h135 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_324); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_326 = 11'h136 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_325); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_327 = 11'h137 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_326); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_328 = 11'h138 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_327); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_329 = 11'h139 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_328); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_330 = 11'h13a == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_329); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_331 = 11'h13b == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_330); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_332 = 11'h13c == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_331); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_333 = 11'h13d == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_332); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_334 = 11'h13e == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_333); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_335 = 11'h13f == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_334); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_336 = 11'h140 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_335); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_337 = 11'h141 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_336); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_338 = 11'h142 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_337); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_339 = 11'h143 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_338); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_340 = 11'h144 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_339); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_341 = 11'h145 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_340); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_342 = 11'h146 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_341); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_343 = 11'h147 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_342); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_344 = 11'h148 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_343); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_345 = 11'h149 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_344); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_346 = 11'h14a == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_345); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_347 = 11'h14b == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_346); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_348 = 11'h14c == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_347); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_349 = 11'h14d == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_348); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_350 = 11'h14e == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_349); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_351 = 11'h14f == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_350); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_352 = 11'h150 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_351); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_353 = 11'h151 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_352); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_354 = 11'h152 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_353); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_355 = 11'h153 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_354); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_356 = 11'h154 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_355); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_357 = 11'h155 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_356); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_358 = 11'h156 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_357); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_359 = 11'h157 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_358); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_360 = 11'h158 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_359); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_361 = 11'h159 == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_360); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_362 = 11'h15a == data2In_0[10:0] ? $signed(5'sh2) : $signed(_GEN_361); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_363 = 11'h15b == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_362); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_364 = 11'h15c == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_363); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_365 = 11'h15d == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_364); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_366 = 11'h15e == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_365); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_367 = 11'h15f == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_366); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_368 = 11'h160 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_367); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_369 = 11'h161 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_368); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_370 = 11'h162 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_369); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_371 = 11'h163 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_370); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_372 = 11'h164 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_371); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_373 = 11'h165 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_372); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_374 = 11'h166 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_373); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_375 = 11'h167 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_374); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_376 = 11'h168 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_375); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_377 = 11'h169 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_376); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_378 = 11'h16a == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_377); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_379 = 11'h16b == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_378); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_380 = 11'h16c == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_379); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_381 = 11'h16d == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_380); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_382 = 11'h16e == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_381); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_383 = 11'h16f == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_382); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_384 = 11'h170 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_383); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_385 = 11'h171 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_384); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_386 = 11'h172 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_385); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_387 = 11'h173 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_386); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_388 = 11'h174 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_387); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_389 = 11'h175 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_388); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_390 = 11'h176 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_389); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_391 = 11'h177 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_390); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_392 = 11'h178 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_391); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_393 = 11'h179 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_392); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_394 = 11'h17a == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_393); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_395 = 11'h17b == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_394); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_396 = 11'h17c == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_395); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_397 = 11'h17d == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_396); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_398 = 11'h17e == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_397); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_399 = 11'h17f == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_398); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_400 = 11'h180 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_399); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_401 = 11'h181 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_400); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_402 = 11'h182 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_401); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_403 = 11'h183 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_402); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_404 = 11'h184 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_403); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_405 = 11'h185 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_404); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_406 = 11'h186 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_405); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_407 = 11'h187 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_406); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_408 = 11'h188 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_407); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_409 = 11'h189 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_408); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_410 = 11'h18a == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_409); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_411 = 11'h18b == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_410); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_412 = 11'h18c == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_411); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_413 = 11'h18d == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_412); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_414 = 11'h18e == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_413); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_415 = 11'h18f == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_414); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_416 = 11'h190 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_415); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_417 = 11'h191 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_416); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_418 = 11'h192 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_417); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_419 = 11'h193 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_418); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_420 = 11'h194 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_419); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_421 = 11'h195 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_420); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_422 = 11'h196 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_421); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_423 = 11'h197 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_422); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_424 = 11'h198 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_423); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_425 = 11'h199 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_424); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_426 = 11'h19a == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_425); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_427 = 11'h19b == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_426); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_428 = 11'h19c == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_427); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_429 = 11'h19d == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_428); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_430 = 11'h19e == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_429); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_431 = 11'h19f == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_430); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_432 = 11'h1a0 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_431); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_433 = 11'h1a1 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_432); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_434 = 11'h1a2 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_433); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_435 = 11'h1a3 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_434); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_436 = 11'h1a4 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_435); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_437 = 11'h1a5 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_436); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_438 = 11'h1a6 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_437); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_439 = 11'h1a7 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_438); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_440 = 11'h1a8 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_439); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_441 = 11'h1a9 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_440); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_442 = 11'h1aa == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_441); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_443 = 11'h1ab == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_442); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_444 = 11'h1ac == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_443); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_445 = 11'h1ad == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_444); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_446 = 11'h1ae == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_445); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_447 = 11'h1af == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_446); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_448 = 11'h1b0 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_447); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_449 = 11'h1b1 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_448); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_450 = 11'h1b2 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_449); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_451 = 11'h1b3 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_450); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_452 = 11'h1b4 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_451); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_453 = 11'h1b5 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_452); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_454 = 11'h1b6 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_453); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_455 = 11'h1b7 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_454); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_456 = 11'h1b8 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_455); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_457 = 11'h1b9 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_456); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_458 = 11'h1ba == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_457); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_459 = 11'h1bb == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_458); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_460 = 11'h1bc == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_459); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_461 = 11'h1bd == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_460); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_462 = 11'h1be == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_461); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_463 = 11'h1bf == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_462); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_464 = 11'h1c0 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_463); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_465 = 11'h1c1 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_464); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_466 = 11'h1c2 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_465); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_467 = 11'h1c3 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_466); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_468 = 11'h1c4 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_467); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_469 = 11'h1c5 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_468); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_470 = 11'h1c6 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_469); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_471 = 11'h1c7 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_470); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_472 = 11'h1c8 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_471); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_473 = 11'h1c9 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_472); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_474 = 11'h1ca == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_473); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_475 = 11'h1cb == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_474); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_476 = 11'h1cc == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_475); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_477 = 11'h1cd == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_476); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_478 = 11'h1ce == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_477); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_479 = 11'h1cf == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_478); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_480 = 11'h1d0 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_479); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_481 = 11'h1d1 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_480); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_482 = 11'h1d2 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_481); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_483 = 11'h1d3 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_482); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_484 = 11'h1d4 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_483); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_485 = 11'h1d5 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_484); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_486 = 11'h1d6 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_485); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_487 = 11'h1d7 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_486); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_488 = 11'h1d8 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_487); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_489 = 11'h1d9 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_488); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_490 = 11'h1da == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_489); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_491 = 11'h1db == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_490); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_492 = 11'h1dc == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_491); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_493 = 11'h1dd == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_492); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_494 = 11'h1de == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_493); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_495 = 11'h1df == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_494); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_496 = 11'h1e0 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_495); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_497 = 11'h1e1 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_496); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_498 = 11'h1e2 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_497); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_499 = 11'h1e3 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_498); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_500 = 11'h1e4 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_499); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_501 = 11'h1e5 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_500); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_502 = 11'h1e6 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_501); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_503 = 11'h1e7 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_502); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_504 = 11'h1e8 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_503); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_505 = 11'h1e9 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_504); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_506 = 11'h1ea == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_505); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_507 = 11'h1eb == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_506); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_508 = 11'h1ec == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_507); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_509 = 11'h1ed == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_508); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_510 = 11'h1ee == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_509); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_511 = 11'h1ef == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_510); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_512 = 11'h1f0 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_511); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_513 = 11'h1f1 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_512); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_514 = 11'h1f2 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_513); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_515 = 11'h1f3 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_514); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_516 = 11'h1f4 == data2In_0[10:0] ? $signed(5'sh3) : $signed(_GEN_515); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_517 = 11'h1f5 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_516); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_518 = 11'h1f6 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_517); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_519 = 11'h1f7 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_518); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_520 = 11'h1f8 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_519); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_521 = 11'h1f9 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_520); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_522 = 11'h1fa == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_521); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_523 = 11'h1fb == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_522); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_524 = 11'h1fc == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_523); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_525 = 11'h1fd == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_524); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_526 = 11'h1fe == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_525); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_527 = 11'h1ff == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_526); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_528 = 11'h200 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_527); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_529 = 11'h201 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_528); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_530 = 11'h202 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_529); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_531 = 11'h203 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_530); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_532 = 11'h204 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_531); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_533 = 11'h205 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_532); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_534 = 11'h206 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_533); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_535 = 11'h207 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_534); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_536 = 11'h208 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_535); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_537 = 11'h209 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_536); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_538 = 11'h20a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_537); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_539 = 11'h20b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_538); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_540 = 11'h20c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_539); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_541 = 11'h20d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_540); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_542 = 11'h20e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_541); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_543 = 11'h20f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_542); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_544 = 11'h210 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_543); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_545 = 11'h211 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_544); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_546 = 11'h212 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_545); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_547 = 11'h213 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_546); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_548 = 11'h214 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_547); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_549 = 11'h215 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_548); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_550 = 11'h216 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_549); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_551 = 11'h217 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_550); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_552 = 11'h218 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_551); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_553 = 11'h219 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_552); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_554 = 11'h21a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_553); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_555 = 11'h21b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_554); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_556 = 11'h21c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_555); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_557 = 11'h21d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_556); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_558 = 11'h21e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_557); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_559 = 11'h21f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_558); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_560 = 11'h220 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_559); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_561 = 11'h221 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_560); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_562 = 11'h222 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_561); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_563 = 11'h223 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_562); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_564 = 11'h224 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_563); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_565 = 11'h225 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_564); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_566 = 11'h226 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_565); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_567 = 11'h227 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_566); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_568 = 11'h228 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_567); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_569 = 11'h229 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_568); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_570 = 11'h22a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_569); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_571 = 11'h22b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_570); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_572 = 11'h22c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_571); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_573 = 11'h22d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_572); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_574 = 11'h22e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_573); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_575 = 11'h22f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_574); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_576 = 11'h230 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_575); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_577 = 11'h231 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_576); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_578 = 11'h232 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_577); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_579 = 11'h233 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_578); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_580 = 11'h234 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_579); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_581 = 11'h235 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_580); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_582 = 11'h236 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_581); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_583 = 11'h237 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_582); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_584 = 11'h238 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_583); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_585 = 11'h239 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_584); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_586 = 11'h23a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_585); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_587 = 11'h23b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_586); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_588 = 11'h23c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_587); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_589 = 11'h23d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_588); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_590 = 11'h23e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_589); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_591 = 11'h23f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_590); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_592 = 11'h240 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_591); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_593 = 11'h241 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_592); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_594 = 11'h242 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_593); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_595 = 11'h243 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_594); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_596 = 11'h244 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_595); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_597 = 11'h245 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_596); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_598 = 11'h246 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_597); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_599 = 11'h247 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_598); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_600 = 11'h248 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_599); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_601 = 11'h249 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_600); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_602 = 11'h24a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_601); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_603 = 11'h24b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_602); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_604 = 11'h24c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_603); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_605 = 11'h24d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_604); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_606 = 11'h24e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_605); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_607 = 11'h24f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_606); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_608 = 11'h250 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_607); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_609 = 11'h251 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_608); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_610 = 11'h252 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_609); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_611 = 11'h253 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_610); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_612 = 11'h254 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_611); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_613 = 11'h255 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_612); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_614 = 11'h256 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_613); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_615 = 11'h257 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_614); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_616 = 11'h258 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_615); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_617 = 11'h259 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_616); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_618 = 11'h25a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_617); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_619 = 11'h25b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_618); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_620 = 11'h25c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_619); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_621 = 11'h25d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_620); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_622 = 11'h25e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_621); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_623 = 11'h25f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_622); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_624 = 11'h260 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_623); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_625 = 11'h261 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_624); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_626 = 11'h262 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_625); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_627 = 11'h263 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_626); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_628 = 11'h264 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_627); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_629 = 11'h265 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_628); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_630 = 11'h266 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_629); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_631 = 11'h267 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_630); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_632 = 11'h268 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_631); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_633 = 11'h269 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_632); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_634 = 11'h26a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_633); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_635 = 11'h26b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_634); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_636 = 11'h26c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_635); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_637 = 11'h26d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_636); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_638 = 11'h26e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_637); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_639 = 11'h26f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_638); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_640 = 11'h270 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_639); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_641 = 11'h271 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_640); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_642 = 11'h272 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_641); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_643 = 11'h273 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_642); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_644 = 11'h274 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_643); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_645 = 11'h275 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_644); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_646 = 11'h276 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_645); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_647 = 11'h277 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_646); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_648 = 11'h278 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_647); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_649 = 11'h279 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_648); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_650 = 11'h27a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_649); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_651 = 11'h27b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_650); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_652 = 11'h27c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_651); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_653 = 11'h27d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_652); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_654 = 11'h27e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_653); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_655 = 11'h27f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_654); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_656 = 11'h280 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_655); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_657 = 11'h281 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_656); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_658 = 11'h282 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_657); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_659 = 11'h283 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_658); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_660 = 11'h284 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_659); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_661 = 11'h285 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_660); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_662 = 11'h286 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_661); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_663 = 11'h287 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_662); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_664 = 11'h288 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_663); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_665 = 11'h289 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_664); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_666 = 11'h28a == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_665); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_667 = 11'h28b == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_666); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_668 = 11'h28c == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_667); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_669 = 11'h28d == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_668); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_670 = 11'h28e == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_669); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_671 = 11'h28f == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_670); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_672 = 11'h290 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_671); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_673 = 11'h291 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_672); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_674 = 11'h292 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_673); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_675 = 11'h293 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_674); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_676 = 11'h294 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_675); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_677 = 11'h295 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_676); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_678 = 11'h296 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_677); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_679 = 11'h297 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_678); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_680 = 11'h298 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_679); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_681 = 11'h299 == data2In_0[10:0] ? $signed(5'sh4) : $signed(_GEN_680); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_682 = 11'h29a == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_681); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_683 = 11'h29b == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_682); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_684 = 11'h29c == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_683); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_685 = 11'h29d == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_684); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_686 = 11'h29e == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_685); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_687 = 11'h29f == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_686); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_688 = 11'h2a0 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_687); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_689 = 11'h2a1 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_688); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_690 = 11'h2a2 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_689); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_691 = 11'h2a3 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_690); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_692 = 11'h2a4 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_691); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_693 = 11'h2a5 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_692); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_694 = 11'h2a6 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_693); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_695 = 11'h2a7 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_694); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_696 = 11'h2a8 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_695); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_697 = 11'h2a9 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_696); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_698 = 11'h2aa == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_697); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_699 = 11'h2ab == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_698); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_700 = 11'h2ac == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_699); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_701 = 11'h2ad == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_700); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_702 = 11'h2ae == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_701); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_703 = 11'h2af == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_702); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_704 = 11'h2b0 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_703); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_705 = 11'h2b1 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_704); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_706 = 11'h2b2 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_705); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_707 = 11'h2b3 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_706); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_708 = 11'h2b4 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_707); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_709 = 11'h2b5 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_708); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_710 = 11'h2b6 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_709); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_711 = 11'h2b7 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_710); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_712 = 11'h2b8 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_711); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_713 = 11'h2b9 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_712); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_714 = 11'h2ba == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_713); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_715 = 11'h2bb == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_714); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_716 = 11'h2bc == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_715); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_717 = 11'h2bd == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_716); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_718 = 11'h2be == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_717); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_719 = 11'h2bf == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_718); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_720 = 11'h2c0 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_719); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_721 = 11'h2c1 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_720); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_722 = 11'h2c2 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_721); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_723 = 11'h2c3 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_722); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_724 = 11'h2c4 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_723); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_725 = 11'h2c5 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_724); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_726 = 11'h2c6 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_725); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_727 = 11'h2c7 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_726); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_728 = 11'h2c8 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_727); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_729 = 11'h2c9 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_728); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_730 = 11'h2ca == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_729); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_731 = 11'h2cb == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_730); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_732 = 11'h2cc == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_731); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_733 = 11'h2cd == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_732); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_734 = 11'h2ce == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_733); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_735 = 11'h2cf == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_734); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_736 = 11'h2d0 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_735); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_737 = 11'h2d1 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_736); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_738 = 11'h2d2 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_737); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_739 = 11'h2d3 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_738); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_740 = 11'h2d4 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_739); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_741 = 11'h2d5 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_740); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_742 = 11'h2d6 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_741); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_743 = 11'h2d7 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_742); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_744 = 11'h2d8 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_743); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_745 = 11'h2d9 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_744); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_746 = 11'h2da == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_745); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_747 = 11'h2db == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_746); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_748 = 11'h2dc == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_747); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_749 = 11'h2dd == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_748); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_750 = 11'h2de == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_749); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_751 = 11'h2df == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_750); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_752 = 11'h2e0 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_751); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_753 = 11'h2e1 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_752); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_754 = 11'h2e2 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_753); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_755 = 11'h2e3 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_754); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_756 = 11'h2e4 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_755); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_757 = 11'h2e5 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_756); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_758 = 11'h2e6 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_757); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_759 = 11'h2e7 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_758); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_760 = 11'h2e8 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_759); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_761 = 11'h2e9 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_760); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_762 = 11'h2ea == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_761); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_763 = 11'h2eb == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_762); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_764 = 11'h2ec == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_763); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_765 = 11'h2ed == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_764); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_766 = 11'h2ee == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_765); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_767 = 11'h2ef == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_766); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_768 = 11'h2f0 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_767); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_769 = 11'h2f1 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_768); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_770 = 11'h2f2 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_769); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_771 = 11'h2f3 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_770); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_772 = 11'h2f4 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_771); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_773 = 11'h2f5 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_772); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_774 = 11'h2f6 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_773); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_775 = 11'h2f7 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_774); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_776 = 11'h2f8 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_775); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_777 = 11'h2f9 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_776); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_778 = 11'h2fa == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_777); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_779 = 11'h2fb == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_778); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_780 = 11'h2fc == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_779); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_781 = 11'h2fd == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_780); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_782 = 11'h2fe == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_781); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_783 = 11'h2ff == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_782); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_784 = 11'h300 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_783); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_785 = 11'h301 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_784); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_786 = 11'h302 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_785); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_787 = 11'h303 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_786); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_788 = 11'h304 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_787); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_789 = 11'h305 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_788); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_790 = 11'h306 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_789); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_791 = 11'h307 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_790); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_792 = 11'h308 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_791); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_793 = 11'h309 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_792); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_794 = 11'h30a == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_793); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_795 = 11'h30b == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_794); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_796 = 11'h30c == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_795); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_797 = 11'h30d == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_796); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_798 = 11'h30e == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_797); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_799 = 11'h30f == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_798); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_800 = 11'h310 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_799); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_801 = 11'h311 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_800); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_802 = 11'h312 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_801); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_803 = 11'h313 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_802); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_804 = 11'h314 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_803); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_805 = 11'h315 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_804); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_806 = 11'h316 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_805); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_807 = 11'h317 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_806); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_808 = 11'h318 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_807); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_809 = 11'h319 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_808); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_810 = 11'h31a == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_809); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_811 = 11'h31b == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_810); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_812 = 11'h31c == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_811); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_813 = 11'h31d == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_812); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_814 = 11'h31e == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_813); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_815 = 11'h31f == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_814); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_816 = 11'h320 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_815); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_817 = 11'h321 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_816); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_818 = 11'h322 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_817); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_819 = 11'h323 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_818); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_820 = 11'h324 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_819); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_821 = 11'h325 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_820); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_822 = 11'h326 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_821); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_823 = 11'h327 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_822); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_824 = 11'h328 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_823); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_825 = 11'h329 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_824); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_826 = 11'h32a == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_825); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_827 = 11'h32b == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_826); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_828 = 11'h32c == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_827); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_829 = 11'h32d == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_828); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_830 = 11'h32e == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_829); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_831 = 11'h32f == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_830); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_832 = 11'h330 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_831); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_833 = 11'h331 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_832); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_834 = 11'h332 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_833); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_835 = 11'h333 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_834); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_836 = 11'h334 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_835); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_837 = 11'h335 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_836); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_838 = 11'h336 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_837); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_839 = 11'h337 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_838); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_840 = 11'h338 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_839); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_841 = 11'h339 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_840); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_842 = 11'h33a == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_841); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_843 = 11'h33b == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_842); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_844 = 11'h33c == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_843); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_845 = 11'h33d == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_844); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_846 = 11'h33e == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_845); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_847 = 11'h33f == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_846); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_848 = 11'h340 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_847); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_849 = 11'h341 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_848); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_850 = 11'h342 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_849); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_851 = 11'h343 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_850); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_852 = 11'h344 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_851); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_853 = 11'h345 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_852); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_854 = 11'h346 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_853); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_855 = 11'h347 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_854); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_856 = 11'h348 == data2In_0[10:0] ? $signed(5'sh5) : $signed(_GEN_855); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_857 = 11'h349 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_856); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_858 = 11'h34a == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_857); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_859 = 11'h34b == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_858); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_860 = 11'h34c == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_859); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_861 = 11'h34d == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_860); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_862 = 11'h34e == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_861); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_863 = 11'h34f == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_862); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_864 = 11'h350 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_863); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_865 = 11'h351 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_864); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_866 = 11'h352 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_865); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_867 = 11'h353 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_866); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_868 = 11'h354 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_867); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_869 = 11'h355 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_868); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_870 = 11'h356 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_869); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_871 = 11'h357 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_870); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_872 = 11'h358 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_871); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_873 = 11'h359 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_872); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_874 = 11'h35a == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_873); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_875 = 11'h35b == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_874); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_876 = 11'h35c == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_875); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_877 = 11'h35d == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_876); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_878 = 11'h35e == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_877); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_879 = 11'h35f == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_878); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_880 = 11'h360 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_879); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_881 = 11'h361 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_880); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_882 = 11'h362 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_881); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_883 = 11'h363 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_882); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_884 = 11'h364 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_883); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_885 = 11'h365 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_884); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_886 = 11'h366 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_885); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_887 = 11'h367 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_886); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_888 = 11'h368 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_887); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_889 = 11'h369 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_888); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_890 = 11'h36a == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_889); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_891 = 11'h36b == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_890); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_892 = 11'h36c == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_891); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_893 = 11'h36d == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_892); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_894 = 11'h36e == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_893); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_895 = 11'h36f == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_894); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_896 = 11'h370 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_895); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_897 = 11'h371 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_896); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_898 = 11'h372 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_897); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_899 = 11'h373 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_898); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_900 = 11'h374 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_899); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_901 = 11'h375 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_900); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_902 = 11'h376 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_901); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_903 = 11'h377 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_902); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_904 = 11'h378 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_903); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_905 = 11'h379 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_904); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_906 = 11'h37a == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_905); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_907 = 11'h37b == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_906); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_908 = 11'h37c == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_907); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_909 = 11'h37d == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_908); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_910 = 11'h37e == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_909); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_911 = 11'h37f == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_910); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_912 = 11'h380 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_911); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_913 = 11'h381 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_912); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_914 = 11'h382 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_913); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_915 = 11'h383 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_914); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_916 = 11'h384 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_915); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_917 = 11'h385 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_916); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_918 = 11'h386 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_917); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_919 = 11'h387 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_918); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_920 = 11'h388 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_919); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_921 = 11'h389 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_920); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_922 = 11'h38a == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_921); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_923 = 11'h38b == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_922); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_924 = 11'h38c == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_923); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_925 = 11'h38d == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_924); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_926 = 11'h38e == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_925); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_927 = 11'h38f == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_926); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_928 = 11'h390 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_927); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_929 = 11'h391 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_928); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_930 = 11'h392 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_929); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_931 = 11'h393 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_930); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_932 = 11'h394 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_931); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_933 = 11'h395 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_932); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_934 = 11'h396 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_933); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_935 = 11'h397 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_934); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_936 = 11'h398 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_935); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_937 = 11'h399 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_936); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_938 = 11'h39a == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_937); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_939 = 11'h39b == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_938); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_940 = 11'h39c == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_939); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_941 = 11'h39d == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_940); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_942 = 11'h39e == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_941); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_943 = 11'h39f == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_942); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_944 = 11'h3a0 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_943); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_945 = 11'h3a1 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_944); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_946 = 11'h3a2 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_945); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_947 = 11'h3a3 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_946); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_948 = 11'h3a4 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_947); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_949 = 11'h3a5 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_948); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_950 = 11'h3a6 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_949); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_951 = 11'h3a7 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_950); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_952 = 11'h3a8 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_951); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_953 = 11'h3a9 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_952); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_954 = 11'h3aa == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_953); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_955 = 11'h3ab == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_954); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_956 = 11'h3ac == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_955); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_957 = 11'h3ad == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_956); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_958 = 11'h3ae == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_957); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_959 = 11'h3af == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_958); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_960 = 11'h3b0 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_959); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_961 = 11'h3b1 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_960); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_962 = 11'h3b2 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_961); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_963 = 11'h3b3 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_962); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_964 = 11'h3b4 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_963); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_965 = 11'h3b5 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_964); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_966 = 11'h3b6 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_965); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_967 = 11'h3b7 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_966); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_968 = 11'h3b8 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_967); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_969 = 11'h3b9 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_968); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_970 = 11'h3ba == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_969); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_971 = 11'h3bb == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_970); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_972 = 11'h3bc == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_971); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_973 = 11'h3bd == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_972); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_974 = 11'h3be == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_973); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_975 = 11'h3bf == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_974); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_976 = 11'h3c0 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_975); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_977 = 11'h3c1 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_976); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_978 = 11'h3c2 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_977); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_979 = 11'h3c3 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_978); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_980 = 11'h3c4 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_979); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_981 = 11'h3c5 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_980); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_982 = 11'h3c6 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_981); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_983 = 11'h3c7 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_982); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_984 = 11'h3c8 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_983); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_985 = 11'h3c9 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_984); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_986 = 11'h3ca == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_985); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_987 = 11'h3cb == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_986); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_988 = 11'h3cc == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_987); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_989 = 11'h3cd == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_988); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_990 = 11'h3ce == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_989); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_991 = 11'h3cf == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_990); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_992 = 11'h3d0 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_991); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_993 = 11'h3d1 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_992); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_994 = 11'h3d2 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_993); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_995 = 11'h3d3 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_994); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_996 = 11'h3d4 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_995); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_997 = 11'h3d5 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_996); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_998 = 11'h3d6 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_997); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_999 = 11'h3d7 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_998); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1000 = 11'h3d8 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_999); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1001 = 11'h3d9 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1000); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1002 = 11'h3da == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1001); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1003 = 11'h3db == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1002); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1004 = 11'h3dc == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1003); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1005 = 11'h3dd == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1004); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1006 = 11'h3de == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1005); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1007 = 11'h3df == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1006); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1008 = 11'h3e0 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1007); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1009 = 11'h3e1 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1008); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1010 = 11'h3e2 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1009); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1011 = 11'h3e3 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1010); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1012 = 11'h3e4 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1011); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1013 = 11'h3e5 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1012); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1014 = 11'h3e6 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1013); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1015 = 11'h3e7 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1014); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1016 = 11'h3e8 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1015); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1017 = 11'h3e9 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1016); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1018 = 11'h3ea == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1017); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1019 = 11'h3eb == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1018); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1020 = 11'h3ec == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1019); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1021 = 11'h3ed == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1020); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1022 = 11'h3ee == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1021); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1023 = 11'h3ef == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1022); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1024 = 11'h3f0 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1023); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1025 = 11'h3f1 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1024); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1026 = 11'h3f2 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1025); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1027 = 11'h3f3 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1026); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1028 = 11'h3f4 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1027); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1029 = 11'h3f5 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1028); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1030 = 11'h3f6 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1029); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1031 = 11'h3f7 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1030); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1032 = 11'h3f8 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1031); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1033 = 11'h3f9 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1032); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1034 = 11'h3fa == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1033); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1035 = 11'h3fb == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1034); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1036 = 11'h3fc == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1035); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1037 = 11'h3fd == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1036); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1038 = 11'h3fe == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1037); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1039 = 11'h3ff == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1038); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1040 = 11'h400 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1039); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1041 = 11'h401 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1040); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1042 = 11'h402 == data2In_0[10:0] ? $signed(5'sh6) : $signed(_GEN_1041); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1043 = 11'h403 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1042); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1044 = 11'h404 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1043); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1045 = 11'h405 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1044); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1046 = 11'h406 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1045); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1047 = 11'h407 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1046); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1048 = 11'h408 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1047); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1049 = 11'h409 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1048); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1050 = 11'h40a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1049); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1051 = 11'h40b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1050); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1052 = 11'h40c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1051); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1053 = 11'h40d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1052); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1054 = 11'h40e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1053); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1055 = 11'h40f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1054); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1056 = 11'h410 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1055); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1057 = 11'h411 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1056); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1058 = 11'h412 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1057); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1059 = 11'h413 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1058); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1060 = 11'h414 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1059); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1061 = 11'h415 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1060); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1062 = 11'h416 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1061); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1063 = 11'h417 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1062); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1064 = 11'h418 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1063); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1065 = 11'h419 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1064); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1066 = 11'h41a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1065); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1067 = 11'h41b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1066); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1068 = 11'h41c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1067); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1069 = 11'h41d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1068); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1070 = 11'h41e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1069); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1071 = 11'h41f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1070); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1072 = 11'h420 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1071); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1073 = 11'h421 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1072); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1074 = 11'h422 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1073); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1075 = 11'h423 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1074); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1076 = 11'h424 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1075); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1077 = 11'h425 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1076); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1078 = 11'h426 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1077); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1079 = 11'h427 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1078); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1080 = 11'h428 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1079); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1081 = 11'h429 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1080); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1082 = 11'h42a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1081); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1083 = 11'h42b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1082); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1084 = 11'h42c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1083); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1085 = 11'h42d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1084); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1086 = 11'h42e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1085); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1087 = 11'h42f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1086); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1088 = 11'h430 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1087); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1089 = 11'h431 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1088); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1090 = 11'h432 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1089); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1091 = 11'h433 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1090); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1092 = 11'h434 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1091); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1093 = 11'h435 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1092); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1094 = 11'h436 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1093); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1095 = 11'h437 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1094); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1096 = 11'h438 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1095); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1097 = 11'h439 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1096); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1098 = 11'h43a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1097); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1099 = 11'h43b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1098); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1100 = 11'h43c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1099); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1101 = 11'h43d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1100); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1102 = 11'h43e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1101); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1103 = 11'h43f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1102); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1104 = 11'h440 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1103); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1105 = 11'h441 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1104); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1106 = 11'h442 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1105); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1107 = 11'h443 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1106); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1108 = 11'h444 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1107); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1109 = 11'h445 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1108); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1110 = 11'h446 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1109); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1111 = 11'h447 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1110); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1112 = 11'h448 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1111); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1113 = 11'h449 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1112); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1114 = 11'h44a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1113); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1115 = 11'h44b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1114); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1116 = 11'h44c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1115); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1117 = 11'h44d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1116); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1118 = 11'h44e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1117); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1119 = 11'h44f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1118); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1120 = 11'h450 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1119); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1121 = 11'h451 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1120); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1122 = 11'h452 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1121); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1123 = 11'h453 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1122); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1124 = 11'h454 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1123); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1125 = 11'h455 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1124); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1126 = 11'h456 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1125); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1127 = 11'h457 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1126); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1128 = 11'h458 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1127); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1129 = 11'h459 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1128); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1130 = 11'h45a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1129); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1131 = 11'h45b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1130); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1132 = 11'h45c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1131); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1133 = 11'h45d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1132); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1134 = 11'h45e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1133); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1135 = 11'h45f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1134); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1136 = 11'h460 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1135); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1137 = 11'h461 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1136); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1138 = 11'h462 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1137); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1139 = 11'h463 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1138); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1140 = 11'h464 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1139); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1141 = 11'h465 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1140); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1142 = 11'h466 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1141); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1143 = 11'h467 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1142); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1144 = 11'h468 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1143); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1145 = 11'h469 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1144); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1146 = 11'h46a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1145); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1147 = 11'h46b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1146); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1148 = 11'h46c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1147); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1149 = 11'h46d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1148); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1150 = 11'h46e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1149); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1151 = 11'h46f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1150); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1152 = 11'h470 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1151); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1153 = 11'h471 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1152); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1154 = 11'h472 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1153); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1155 = 11'h473 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1154); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1156 = 11'h474 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1155); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1157 = 11'h475 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1156); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1158 = 11'h476 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1157); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1159 = 11'h477 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1158); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1160 = 11'h478 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1159); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1161 = 11'h479 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1160); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1162 = 11'h47a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1161); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1163 = 11'h47b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1162); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1164 = 11'h47c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1163); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1165 = 11'h47d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1164); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1166 = 11'h47e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1165); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1167 = 11'h47f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1166); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1168 = 11'h480 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1167); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1169 = 11'h481 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1168); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1170 = 11'h482 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1169); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1171 = 11'h483 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1170); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1172 = 11'h484 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1171); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1173 = 11'h485 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1172); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1174 = 11'h486 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1173); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1175 = 11'h487 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1174); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1176 = 11'h488 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1175); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1177 = 11'h489 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1176); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1178 = 11'h48a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1177); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1179 = 11'h48b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1178); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1180 = 11'h48c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1179); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1181 = 11'h48d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1180); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1182 = 11'h48e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1181); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1183 = 11'h48f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1182); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1184 = 11'h490 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1183); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1185 = 11'h491 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1184); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1186 = 11'h492 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1185); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1187 = 11'h493 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1186); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1188 = 11'h494 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1187); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1189 = 11'h495 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1188); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1190 = 11'h496 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1189); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1191 = 11'h497 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1190); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1192 = 11'h498 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1191); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1193 = 11'h499 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1192); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1194 = 11'h49a == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1193); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1195 = 11'h49b == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1194); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1196 = 11'h49c == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1195); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1197 = 11'h49d == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1196); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1198 = 11'h49e == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1197); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1199 = 11'h49f == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1198); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1200 = 11'h4a0 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1199); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1201 = 11'h4a1 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1200); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1202 = 11'h4a2 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1201); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1203 = 11'h4a3 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1202); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1204 = 11'h4a4 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1203); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1205 = 11'h4a5 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1204); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1206 = 11'h4a6 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1205); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1207 = 11'h4a7 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1206); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1208 = 11'h4a8 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1207); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1209 = 11'h4a9 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1208); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1210 = 11'h4aa == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1209); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1211 = 11'h4ab == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1210); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1212 = 11'h4ac == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1211); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1213 = 11'h4ad == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1212); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1214 = 11'h4ae == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1213); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1215 = 11'h4af == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1214); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1216 = 11'h4b0 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1215); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1217 = 11'h4b1 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1216); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1218 = 11'h4b2 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1217); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1219 = 11'h4b3 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1218); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1220 = 11'h4b4 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1219); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1221 = 11'h4b5 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1220); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1222 = 11'h4b6 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1221); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1223 = 11'h4b7 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1222); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1224 = 11'h4b8 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1223); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1225 = 11'h4b9 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1224); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1226 = 11'h4ba == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1225); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1227 = 11'h4bb == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1226); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1228 = 11'h4bc == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1227); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1229 = 11'h4bd == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1228); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1230 = 11'h4be == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1229); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1231 = 11'h4bf == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1230); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1232 = 11'h4c0 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1231); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1233 = 11'h4c1 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1232); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1234 = 11'h4c2 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1233); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1235 = 11'h4c3 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1234); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1236 = 11'h4c4 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1235); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1237 = 11'h4c5 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1236); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1238 = 11'h4c6 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1237); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1239 = 11'h4c7 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1238); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1240 = 11'h4c8 == data2In_0[10:0] ? $signed(5'sh7) : $signed(_GEN_1239); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1241 = 11'h4c9 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1240); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1242 = 11'h4ca == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1241); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1243 = 11'h4cb == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1242); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1244 = 11'h4cc == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1243); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1245 = 11'h4cd == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1244); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1246 = 11'h4ce == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1245); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1247 = 11'h4cf == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1246); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1248 = 11'h4d0 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1247); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1249 = 11'h4d1 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1248); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1250 = 11'h4d2 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1249); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1251 = 11'h4d3 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1250); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1252 = 11'h4d4 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1251); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1253 = 11'h4d5 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1252); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1254 = 11'h4d6 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1253); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1255 = 11'h4d7 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1254); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1256 = 11'h4d8 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1255); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1257 = 11'h4d9 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1256); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1258 = 11'h4da == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1257); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1259 = 11'h4db == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1258); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1260 = 11'h4dc == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1259); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1261 = 11'h4dd == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1260); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1262 = 11'h4de == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1261); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1263 = 11'h4df == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1262); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1264 = 11'h4e0 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1263); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1265 = 11'h4e1 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1264); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1266 = 11'h4e2 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1265); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1267 = 11'h4e3 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1266); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1268 = 11'h4e4 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1267); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1269 = 11'h4e5 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1268); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1270 = 11'h4e6 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1269); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1271 = 11'h4e7 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1270); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1272 = 11'h4e8 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1271); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1273 = 11'h4e9 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1272); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1274 = 11'h4ea == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1273); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1275 = 11'h4eb == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1274); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1276 = 11'h4ec == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1275); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1277 = 11'h4ed == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1276); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1278 = 11'h4ee == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1277); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1279 = 11'h4ef == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1278); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1280 = 11'h4f0 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1279); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1281 = 11'h4f1 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1280); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1282 = 11'h4f2 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1281); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1283 = 11'h4f3 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1282); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1284 = 11'h4f4 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1283); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1285 = 11'h4f5 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1284); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1286 = 11'h4f6 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1285); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1287 = 11'h4f7 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1286); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1288 = 11'h4f8 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1287); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1289 = 11'h4f9 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1288); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1290 = 11'h4fa == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1289); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1291 = 11'h4fb == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1290); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1292 = 11'h4fc == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1291); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1293 = 11'h4fd == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1292); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1294 = 11'h4fe == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1293); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1295 = 11'h4ff == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1294); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1296 = 11'h500 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1295); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1297 = 11'h501 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1296); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1298 = 11'h502 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1297); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1299 = 11'h503 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1298); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1300 = 11'h504 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1299); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1301 = 11'h505 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1300); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1302 = 11'h506 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1301); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1303 = 11'h507 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1302); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1304 = 11'h508 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1303); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1305 = 11'h509 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1304); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1306 = 11'h50a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1305); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1307 = 11'h50b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1306); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1308 = 11'h50c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1307); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1309 = 11'h50d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1308); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1310 = 11'h50e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1309); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1311 = 11'h50f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1310); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1312 = 11'h510 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1311); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1313 = 11'h511 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1312); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1314 = 11'h512 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1313); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1315 = 11'h513 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1314); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1316 = 11'h514 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1315); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1317 = 11'h515 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1316); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1318 = 11'h516 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1317); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1319 = 11'h517 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1318); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1320 = 11'h518 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1319); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1321 = 11'h519 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1320); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1322 = 11'h51a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1321); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1323 = 11'h51b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1322); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1324 = 11'h51c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1323); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1325 = 11'h51d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1324); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1326 = 11'h51e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1325); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1327 = 11'h51f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1326); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1328 = 11'h520 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1327); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1329 = 11'h521 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1328); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1330 = 11'h522 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1329); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1331 = 11'h523 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1330); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1332 = 11'h524 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1331); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1333 = 11'h525 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1332); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1334 = 11'h526 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1333); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1335 = 11'h527 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1334); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1336 = 11'h528 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1335); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1337 = 11'h529 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1336); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1338 = 11'h52a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1337); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1339 = 11'h52b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1338); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1340 = 11'h52c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1339); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1341 = 11'h52d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1340); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1342 = 11'h52e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1341); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1343 = 11'h52f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1342); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1344 = 11'h530 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1343); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1345 = 11'h531 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1344); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1346 = 11'h532 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1345); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1347 = 11'h533 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1346); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1348 = 11'h534 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1347); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1349 = 11'h535 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1348); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1350 = 11'h536 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1349); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1351 = 11'h537 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1350); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1352 = 11'h538 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1351); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1353 = 11'h539 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1352); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1354 = 11'h53a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1353); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1355 = 11'h53b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1354); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1356 = 11'h53c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1355); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1357 = 11'h53d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1356); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1358 = 11'h53e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1357); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1359 = 11'h53f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1358); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1360 = 11'h540 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1359); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1361 = 11'h541 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1360); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1362 = 11'h542 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1361); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1363 = 11'h543 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1362); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1364 = 11'h544 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1363); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1365 = 11'h545 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1364); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1366 = 11'h546 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1365); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1367 = 11'h547 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1366); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1368 = 11'h548 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1367); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1369 = 11'h549 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1368); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1370 = 11'h54a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1369); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1371 = 11'h54b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1370); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1372 = 11'h54c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1371); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1373 = 11'h54d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1372); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1374 = 11'h54e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1373); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1375 = 11'h54f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1374); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1376 = 11'h550 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1375); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1377 = 11'h551 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1376); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1378 = 11'h552 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1377); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1379 = 11'h553 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1378); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1380 = 11'h554 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1379); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1381 = 11'h555 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1380); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1382 = 11'h556 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1381); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1383 = 11'h557 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1382); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1384 = 11'h558 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1383); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1385 = 11'h559 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1384); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1386 = 11'h55a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1385); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1387 = 11'h55b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1386); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1388 = 11'h55c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1387); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1389 = 11'h55d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1388); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1390 = 11'h55e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1389); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1391 = 11'h55f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1390); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1392 = 11'h560 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1391); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1393 = 11'h561 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1392); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1394 = 11'h562 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1393); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1395 = 11'h563 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1394); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1396 = 11'h564 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1395); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1397 = 11'h565 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1396); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1398 = 11'h566 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1397); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1399 = 11'h567 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1398); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1400 = 11'h568 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1399); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1401 = 11'h569 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1400); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1402 = 11'h56a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1401); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1403 = 11'h56b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1402); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1404 = 11'h56c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1403); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1405 = 11'h56d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1404); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1406 = 11'h56e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1405); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1407 = 11'h56f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1406); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1408 = 11'h570 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1407); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1409 = 11'h571 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1408); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1410 = 11'h572 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1409); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1411 = 11'h573 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1410); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1412 = 11'h574 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1411); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1413 = 11'h575 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1412); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1414 = 11'h576 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1413); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1415 = 11'h577 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1414); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1416 = 11'h578 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1415); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1417 = 11'h579 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1416); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1418 = 11'h57a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1417); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1419 = 11'h57b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1418); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1420 = 11'h57c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1419); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1421 = 11'h57d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1420); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1422 = 11'h57e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1421); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1423 = 11'h57f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1422); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1424 = 11'h580 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1423); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1425 = 11'h581 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1424); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1426 = 11'h582 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1425); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1427 = 11'h583 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1426); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1428 = 11'h584 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1427); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1429 = 11'h585 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1428); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1430 = 11'h586 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1429); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1431 = 11'h587 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1430); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1432 = 11'h588 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1431); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1433 = 11'h589 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1432); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1434 = 11'h58a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1433); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1435 = 11'h58b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1434); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1436 = 11'h58c == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1435); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1437 = 11'h58d == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1436); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1438 = 11'h58e == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1437); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1439 = 11'h58f == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1438); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1440 = 11'h590 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1439); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1441 = 11'h591 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1440); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1442 = 11'h592 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1441); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1443 = 11'h593 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1442); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1444 = 11'h594 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1443); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1445 = 11'h595 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1444); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1446 = 11'h596 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1445); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1447 = 11'h597 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1446); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1448 = 11'h598 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1447); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1449 = 11'h599 == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1448); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1450 = 11'h59a == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1449); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1451 = 11'h59b == data2In_0[10:0] ? $signed(5'sh8) : $signed(_GEN_1450); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1452 = 11'h59c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1451); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1453 = 11'h59d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1452); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1454 = 11'h59e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1453); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1455 = 11'h59f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1454); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1456 = 11'h5a0 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1455); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1457 = 11'h5a1 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1456); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1458 = 11'h5a2 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1457); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1459 = 11'h5a3 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1458); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1460 = 11'h5a4 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1459); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1461 = 11'h5a5 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1460); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1462 = 11'h5a6 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1461); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1463 = 11'h5a7 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1462); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1464 = 11'h5a8 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1463); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1465 = 11'h5a9 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1464); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1466 = 11'h5aa == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1465); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1467 = 11'h5ab == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1466); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1468 = 11'h5ac == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1467); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1469 = 11'h5ad == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1468); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1470 = 11'h5ae == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1469); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1471 = 11'h5af == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1470); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1472 = 11'h5b0 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1471); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1473 = 11'h5b1 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1472); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1474 = 11'h5b2 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1473); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1475 = 11'h5b3 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1474); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1476 = 11'h5b4 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1475); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1477 = 11'h5b5 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1476); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1478 = 11'h5b6 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1477); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1479 = 11'h5b7 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1478); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1480 = 11'h5b8 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1479); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1481 = 11'h5b9 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1480); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1482 = 11'h5ba == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1481); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1483 = 11'h5bb == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1482); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1484 = 11'h5bc == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1483); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1485 = 11'h5bd == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1484); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1486 = 11'h5be == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1485); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1487 = 11'h5bf == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1486); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1488 = 11'h5c0 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1487); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1489 = 11'h5c1 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1488); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1490 = 11'h5c2 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1489); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1491 = 11'h5c3 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1490); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1492 = 11'h5c4 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1491); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1493 = 11'h5c5 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1492); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1494 = 11'h5c6 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1493); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1495 = 11'h5c7 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1494); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1496 = 11'h5c8 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1495); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1497 = 11'h5c9 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1496); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1498 = 11'h5ca == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1497); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1499 = 11'h5cb == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1498); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1500 = 11'h5cc == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1499); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1501 = 11'h5cd == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1500); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1502 = 11'h5ce == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1501); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1503 = 11'h5cf == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1502); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1504 = 11'h5d0 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1503); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1505 = 11'h5d1 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1504); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1506 = 11'h5d2 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1505); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1507 = 11'h5d3 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1506); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1508 = 11'h5d4 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1507); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1509 = 11'h5d5 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1508); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1510 = 11'h5d6 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1509); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1511 = 11'h5d7 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1510); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1512 = 11'h5d8 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1511); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1513 = 11'h5d9 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1512); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1514 = 11'h5da == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1513); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1515 = 11'h5db == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1514); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1516 = 11'h5dc == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1515); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1517 = 11'h5dd == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1516); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1518 = 11'h5de == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1517); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1519 = 11'h5df == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1518); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1520 = 11'h5e0 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1519); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1521 = 11'h5e1 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1520); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1522 = 11'h5e2 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1521); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1523 = 11'h5e3 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1522); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1524 = 11'h5e4 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1523); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1525 = 11'h5e5 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1524); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1526 = 11'h5e6 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1525); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1527 = 11'h5e7 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1526); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1528 = 11'h5e8 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1527); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1529 = 11'h5e9 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1528); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1530 = 11'h5ea == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1529); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1531 = 11'h5eb == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1530); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1532 = 11'h5ec == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1531); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1533 = 11'h5ed == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1532); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1534 = 11'h5ee == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1533); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1535 = 11'h5ef == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1534); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1536 = 11'h5f0 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1535); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1537 = 11'h5f1 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1536); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1538 = 11'h5f2 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1537); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1539 = 11'h5f3 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1538); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1540 = 11'h5f4 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1539); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1541 = 11'h5f5 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1540); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1542 = 11'h5f6 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1541); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1543 = 11'h5f7 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1542); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1544 = 11'h5f8 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1543); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1545 = 11'h5f9 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1544); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1546 = 11'h5fa == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1545); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1547 = 11'h5fb == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1546); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1548 = 11'h5fc == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1547); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1549 = 11'h5fd == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1548); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1550 = 11'h5fe == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1549); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1551 = 11'h5ff == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1550); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1552 = 11'h600 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1551); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1553 = 11'h601 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1552); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1554 = 11'h602 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1553); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1555 = 11'h603 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1554); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1556 = 11'h604 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1555); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1557 = 11'h605 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1556); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1558 = 11'h606 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1557); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1559 = 11'h607 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1558); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1560 = 11'h608 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1559); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1561 = 11'h609 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1560); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1562 = 11'h60a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1561); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1563 = 11'h60b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1562); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1564 = 11'h60c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1563); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1565 = 11'h60d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1564); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1566 = 11'h60e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1565); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1567 = 11'h60f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1566); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1568 = 11'h610 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1567); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1569 = 11'h611 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1568); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1570 = 11'h612 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1569); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1571 = 11'h613 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1570); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1572 = 11'h614 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1571); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1573 = 11'h615 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1572); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1574 = 11'h616 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1573); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1575 = 11'h617 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1574); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1576 = 11'h618 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1575); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1577 = 11'h619 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1576); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1578 = 11'h61a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1577); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1579 = 11'h61b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1578); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1580 = 11'h61c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1579); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1581 = 11'h61d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1580); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1582 = 11'h61e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1581); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1583 = 11'h61f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1582); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1584 = 11'h620 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1583); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1585 = 11'h621 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1584); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1586 = 11'h622 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1585); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1587 = 11'h623 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1586); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1588 = 11'h624 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1587); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1589 = 11'h625 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1588); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1590 = 11'h626 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1589); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1591 = 11'h627 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1590); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1592 = 11'h628 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1591); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1593 = 11'h629 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1592); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1594 = 11'h62a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1593); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1595 = 11'h62b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1594); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1596 = 11'h62c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1595); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1597 = 11'h62d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1596); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1598 = 11'h62e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1597); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1599 = 11'h62f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1598); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1600 = 11'h630 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1599); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1601 = 11'h631 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1600); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1602 = 11'h632 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1601); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1603 = 11'h633 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1602); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1604 = 11'h634 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1603); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1605 = 11'h635 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1604); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1606 = 11'h636 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1605); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1607 = 11'h637 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1606); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1608 = 11'h638 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1607); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1609 = 11'h639 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1608); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1610 = 11'h63a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1609); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1611 = 11'h63b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1610); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1612 = 11'h63c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1611); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1613 = 11'h63d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1612); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1614 = 11'h63e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1613); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1615 = 11'h63f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1614); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1616 = 11'h640 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1615); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1617 = 11'h641 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1616); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1618 = 11'h642 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1617); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1619 = 11'h643 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1618); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1620 = 11'h644 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1619); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1621 = 11'h645 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1620); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1622 = 11'h646 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1621); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1623 = 11'h647 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1622); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1624 = 11'h648 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1623); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1625 = 11'h649 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1624); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1626 = 11'h64a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1625); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1627 = 11'h64b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1626); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1628 = 11'h64c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1627); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1629 = 11'h64d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1628); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1630 = 11'h64e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1629); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1631 = 11'h64f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1630); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1632 = 11'h650 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1631); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1633 = 11'h651 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1632); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1634 = 11'h652 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1633); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1635 = 11'h653 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1634); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1636 = 11'h654 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1635); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1637 = 11'h655 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1636); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1638 = 11'h656 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1637); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1639 = 11'h657 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1638); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1640 = 11'h658 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1639); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1641 = 11'h659 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1640); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1642 = 11'h65a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1641); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1643 = 11'h65b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1642); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1644 = 11'h65c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1643); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1645 = 11'h65d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1644); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1646 = 11'h65e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1645); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1647 = 11'h65f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1646); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1648 = 11'h660 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1647); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1649 = 11'h661 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1648); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1650 = 11'h662 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1649); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1651 = 11'h663 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1650); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1652 = 11'h664 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1651); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1653 = 11'h665 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1652); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1654 = 11'h666 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1653); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1655 = 11'h667 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1654); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1656 = 11'h668 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1655); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1657 = 11'h669 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1656); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1658 = 11'h66a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1657); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1659 = 11'h66b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1658); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1660 = 11'h66c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1659); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1661 = 11'h66d == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1660); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1662 = 11'h66e == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1661); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1663 = 11'h66f == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1662); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1664 = 11'h670 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1663); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1665 = 11'h671 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1664); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1666 = 11'h672 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1665); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1667 = 11'h673 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1666); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1668 = 11'h674 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1667); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1669 = 11'h675 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1668); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1670 = 11'h676 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1669); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1671 = 11'h677 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1670); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1672 = 11'h678 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1671); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1673 = 11'h679 == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1672); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1674 = 11'h67a == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1673); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1675 = 11'h67b == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1674); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1676 = 11'h67c == data2In_0[10:0] ? $signed(5'sh9) : $signed(_GEN_1675); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1677 = 11'h67d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1676); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1678 = 11'h67e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1677); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1679 = 11'h67f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1678); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1680 = 11'h680 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1679); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1681 = 11'h681 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1680); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1682 = 11'h682 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1681); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1683 = 11'h683 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1682); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1684 = 11'h684 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1683); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1685 = 11'h685 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1684); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1686 = 11'h686 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1685); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1687 = 11'h687 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1686); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1688 = 11'h688 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1687); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1689 = 11'h689 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1688); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1690 = 11'h68a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1689); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1691 = 11'h68b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1690); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1692 = 11'h68c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1691); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1693 = 11'h68d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1692); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1694 = 11'h68e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1693); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1695 = 11'h68f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1694); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1696 = 11'h690 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1695); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1697 = 11'h691 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1696); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1698 = 11'h692 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1697); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1699 = 11'h693 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1698); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1700 = 11'h694 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1699); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1701 = 11'h695 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1700); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1702 = 11'h696 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1701); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1703 = 11'h697 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1702); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1704 = 11'h698 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1703); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1705 = 11'h699 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1704); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1706 = 11'h69a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1705); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1707 = 11'h69b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1706); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1708 = 11'h69c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1707); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1709 = 11'h69d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1708); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1710 = 11'h69e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1709); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1711 = 11'h69f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1710); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1712 = 11'h6a0 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1711); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1713 = 11'h6a1 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1712); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1714 = 11'h6a2 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1713); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1715 = 11'h6a3 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1714); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1716 = 11'h6a4 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1715); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1717 = 11'h6a5 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1716); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1718 = 11'h6a6 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1717); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1719 = 11'h6a7 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1718); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1720 = 11'h6a8 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1719); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1721 = 11'h6a9 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1720); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1722 = 11'h6aa == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1721); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1723 = 11'h6ab == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1722); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1724 = 11'h6ac == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1723); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1725 = 11'h6ad == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1724); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1726 = 11'h6ae == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1725); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1727 = 11'h6af == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1726); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1728 = 11'h6b0 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1727); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1729 = 11'h6b1 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1728); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1730 = 11'h6b2 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1729); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1731 = 11'h6b3 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1730); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1732 = 11'h6b4 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1731); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1733 = 11'h6b5 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1732); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1734 = 11'h6b6 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1733); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1735 = 11'h6b7 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1734); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1736 = 11'h6b8 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1735); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1737 = 11'h6b9 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1736); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1738 = 11'h6ba == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1737); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1739 = 11'h6bb == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1738); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1740 = 11'h6bc == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1739); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1741 = 11'h6bd == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1740); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1742 = 11'h6be == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1741); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1743 = 11'h6bf == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1742); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1744 = 11'h6c0 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1743); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1745 = 11'h6c1 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1744); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1746 = 11'h6c2 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1745); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1747 = 11'h6c3 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1746); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1748 = 11'h6c4 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1747); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1749 = 11'h6c5 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1748); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1750 = 11'h6c6 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1749); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1751 = 11'h6c7 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1750); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1752 = 11'h6c8 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1751); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1753 = 11'h6c9 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1752); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1754 = 11'h6ca == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1753); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1755 = 11'h6cb == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1754); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1756 = 11'h6cc == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1755); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1757 = 11'h6cd == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1756); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1758 = 11'h6ce == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1757); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1759 = 11'h6cf == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1758); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1760 = 11'h6d0 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1759); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1761 = 11'h6d1 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1760); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1762 = 11'h6d2 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1761); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1763 = 11'h6d3 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1762); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1764 = 11'h6d4 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1763); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1765 = 11'h6d5 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1764); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1766 = 11'h6d6 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1765); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1767 = 11'h6d7 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1766); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1768 = 11'h6d8 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1767); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1769 = 11'h6d9 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1768); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1770 = 11'h6da == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1769); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1771 = 11'h6db == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1770); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1772 = 11'h6dc == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1771); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1773 = 11'h6dd == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1772); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1774 = 11'h6de == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1773); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1775 = 11'h6df == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1774); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1776 = 11'h6e0 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1775); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1777 = 11'h6e1 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1776); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1778 = 11'h6e2 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1777); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1779 = 11'h6e3 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1778); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1780 = 11'h6e4 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1779); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1781 = 11'h6e5 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1780); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1782 = 11'h6e6 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1781); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1783 = 11'h6e7 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1782); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1784 = 11'h6e8 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1783); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1785 = 11'h6e9 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1784); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1786 = 11'h6ea == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1785); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1787 = 11'h6eb == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1786); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1788 = 11'h6ec == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1787); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1789 = 11'h6ed == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1788); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1790 = 11'h6ee == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1789); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1791 = 11'h6ef == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1790); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1792 = 11'h6f0 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1791); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1793 = 11'h6f1 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1792); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1794 = 11'h6f2 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1793); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1795 = 11'h6f3 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1794); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1796 = 11'h6f4 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1795); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1797 = 11'h6f5 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1796); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1798 = 11'h6f6 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1797); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1799 = 11'h6f7 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1798); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1800 = 11'h6f8 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1799); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1801 = 11'h6f9 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1800); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1802 = 11'h6fa == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1801); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1803 = 11'h6fb == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1802); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1804 = 11'h6fc == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1803); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1805 = 11'h6fd == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1804); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1806 = 11'h6fe == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1805); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1807 = 11'h6ff == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1806); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1808 = 11'h700 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1807); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1809 = 11'h701 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1808); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1810 = 11'h702 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1809); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1811 = 11'h703 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1810); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1812 = 11'h704 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1811); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1813 = 11'h705 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1812); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1814 = 11'h706 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1813); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1815 = 11'h707 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1814); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1816 = 11'h708 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1815); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1817 = 11'h709 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1816); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1818 = 11'h70a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1817); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1819 = 11'h70b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1818); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1820 = 11'h70c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1819); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1821 = 11'h70d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1820); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1822 = 11'h70e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1821); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1823 = 11'h70f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1822); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1824 = 11'h710 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1823); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1825 = 11'h711 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1824); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1826 = 11'h712 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1825); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1827 = 11'h713 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1826); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1828 = 11'h714 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1827); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1829 = 11'h715 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1828); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1830 = 11'h716 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1829); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1831 = 11'h717 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1830); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1832 = 11'h718 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1831); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1833 = 11'h719 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1832); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1834 = 11'h71a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1833); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1835 = 11'h71b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1834); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1836 = 11'h71c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1835); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1837 = 11'h71d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1836); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1838 = 11'h71e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1837); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1839 = 11'h71f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1838); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1840 = 11'h720 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1839); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1841 = 11'h721 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1840); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1842 = 11'h722 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1841); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1843 = 11'h723 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1842); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1844 = 11'h724 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1843); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1845 = 11'h725 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1844); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1846 = 11'h726 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1845); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1847 = 11'h727 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1846); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1848 = 11'h728 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1847); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1849 = 11'h729 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1848); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1850 = 11'h72a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1849); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1851 = 11'h72b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1850); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1852 = 11'h72c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1851); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1853 = 11'h72d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1852); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1854 = 11'h72e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1853); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1855 = 11'h72f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1854); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1856 = 11'h730 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1855); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1857 = 11'h731 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1856); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1858 = 11'h732 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1857); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1859 = 11'h733 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1858); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1860 = 11'h734 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1859); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1861 = 11'h735 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1860); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1862 = 11'h736 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1861); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1863 = 11'h737 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1862); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1864 = 11'h738 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1863); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1865 = 11'h739 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1864); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1866 = 11'h73a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1865); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1867 = 11'h73b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1866); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1868 = 11'h73c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1867); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1869 = 11'h73d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1868); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1870 = 11'h73e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1869); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1871 = 11'h73f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1870); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1872 = 11'h740 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1871); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1873 = 11'h741 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1872); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1874 = 11'h742 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1873); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1875 = 11'h743 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1874); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1876 = 11'h744 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1875); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1877 = 11'h745 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1876); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1878 = 11'h746 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1877); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1879 = 11'h747 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1878); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1880 = 11'h748 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1879); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1881 = 11'h749 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1880); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1882 = 11'h74a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1881); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1883 = 11'h74b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1882); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1884 = 11'h74c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1883); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1885 = 11'h74d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1884); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1886 = 11'h74e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1885); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1887 = 11'h74f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1886); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1888 = 11'h750 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1887); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1889 = 11'h751 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1888); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1890 = 11'h752 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1889); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1891 = 11'h753 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1890); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1892 = 11'h754 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1891); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1893 = 11'h755 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1892); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1894 = 11'h756 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1893); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1895 = 11'h757 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1894); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1896 = 11'h758 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1895); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1897 = 11'h759 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1896); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1898 = 11'h75a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1897); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1899 = 11'h75b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1898); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1900 = 11'h75c == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1899); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1901 = 11'h75d == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1900); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1902 = 11'h75e == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1901); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1903 = 11'h75f == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1902); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1904 = 11'h760 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1903); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1905 = 11'h761 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1904); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1906 = 11'h762 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1905); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1907 = 11'h763 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1906); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1908 = 11'h764 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1907); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1909 = 11'h765 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1908); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1910 = 11'h766 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1909); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1911 = 11'h767 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1910); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1912 = 11'h768 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1911); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1913 = 11'h769 == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1912); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1914 = 11'h76a == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1913); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1915 = 11'h76b == data2In_0[10:0] ? $signed(5'sha) : $signed(_GEN_1914); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1916 = 11'h76c == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1915); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1917 = 11'h76d == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1916); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1918 = 11'h76e == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1917); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1919 = 11'h76f == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1918); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1920 = 11'h770 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1919); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1921 = 11'h771 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1920); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1922 = 11'h772 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1921); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1923 = 11'h773 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1922); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1924 = 11'h774 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1923); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1925 = 11'h775 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1924); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1926 = 11'h776 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1925); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1927 = 11'h777 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1926); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1928 = 11'h778 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1927); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1929 = 11'h779 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1928); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1930 = 11'h77a == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1929); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1931 = 11'h77b == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1930); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1932 = 11'h77c == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1931); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1933 = 11'h77d == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1932); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1934 = 11'h77e == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1933); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1935 = 11'h77f == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1934); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1936 = 11'h780 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1935); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1937 = 11'h781 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1936); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1938 = 11'h782 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1937); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1939 = 11'h783 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1938); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1940 = 11'h784 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1939); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1941 = 11'h785 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1940); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1942 = 11'h786 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1941); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1943 = 11'h787 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1942); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1944 = 11'h788 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1943); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1945 = 11'h789 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1944); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1946 = 11'h78a == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1945); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1947 = 11'h78b == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1946); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1948 = 11'h78c == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1947); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1949 = 11'h78d == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1948); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1950 = 11'h78e == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1949); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1951 = 11'h78f == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1950); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1952 = 11'h790 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1951); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1953 = 11'h791 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1952); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1954 = 11'h792 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1953); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1955 = 11'h793 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1954); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1956 = 11'h794 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1955); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1957 = 11'h795 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1956); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1958 = 11'h796 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1957); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1959 = 11'h797 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1958); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1960 = 11'h798 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1959); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1961 = 11'h799 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1960); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1962 = 11'h79a == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1961); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1963 = 11'h79b == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1962); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1964 = 11'h79c == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1963); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1965 = 11'h79d == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1964); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1966 = 11'h79e == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1965); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1967 = 11'h79f == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1966); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1968 = 11'h7a0 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1967); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1969 = 11'h7a1 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1968); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1970 = 11'h7a2 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1969); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1971 = 11'h7a3 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1970); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1972 = 11'h7a4 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1971); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1973 = 11'h7a5 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1972); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1974 = 11'h7a6 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1973); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1975 = 11'h7a7 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1974); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1976 = 11'h7a8 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1975); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1977 = 11'h7a9 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1976); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1978 = 11'h7aa == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1977); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1979 = 11'h7ab == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1978); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1980 = 11'h7ac == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1979); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1981 = 11'h7ad == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1980); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1982 = 11'h7ae == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1981); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1983 = 11'h7af == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1982); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1984 = 11'h7b0 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1983); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1985 = 11'h7b1 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1984); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1986 = 11'h7b2 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1985); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1987 = 11'h7b3 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1986); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1988 = 11'h7b4 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1987); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1989 = 11'h7b5 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1988); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1990 = 11'h7b6 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1989); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1991 = 11'h7b7 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1990); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1992 = 11'h7b8 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1991); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1993 = 11'h7b9 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1992); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1994 = 11'h7ba == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1993); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1995 = 11'h7bb == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1994); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1996 = 11'h7bc == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1995); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1997 = 11'h7bd == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1996); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1998 = 11'h7be == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1997); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_1999 = 11'h7bf == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1998); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2000 = 11'h7c0 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_1999); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2001 = 11'h7c1 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2000); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2002 = 11'h7c2 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2001); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2003 = 11'h7c3 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2002); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2004 = 11'h7c4 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2003); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2005 = 11'h7c5 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2004); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2006 = 11'h7c6 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2005); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2007 = 11'h7c7 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2006); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2008 = 11'h7c8 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2007); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2009 = 11'h7c9 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2008); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2010 = 11'h7ca == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2009); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2011 = 11'h7cb == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2010); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2012 = 11'h7cc == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2011); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2013 = 11'h7cd == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2012); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2014 = 11'h7ce == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2013); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2015 = 11'h7cf == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2014); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2016 = 11'h7d0 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2015); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2017 = 11'h7d1 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2016); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2018 = 11'h7d2 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2017); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2019 = 11'h7d3 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2018); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2020 = 11'h7d4 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2019); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2021 = 11'h7d5 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2020); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2022 = 11'h7d6 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2021); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2023 = 11'h7d7 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2022); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2024 = 11'h7d8 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2023); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2025 = 11'h7d9 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2024); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2026 = 11'h7da == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2025); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2027 = 11'h7db == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2026); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2028 = 11'h7dc == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2027); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2029 = 11'h7dd == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2028); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2030 = 11'h7de == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2029); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2031 = 11'h7df == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2030); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2032 = 11'h7e0 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2031); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2033 = 11'h7e1 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2032); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2034 = 11'h7e2 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2033); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2035 = 11'h7e3 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2034); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2036 = 11'h7e4 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2035); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2037 = 11'h7e5 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2036); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2038 = 11'h7e6 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2037); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2039 = 11'h7e7 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2038); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2040 = 11'h7e8 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2039); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2041 = 11'h7e9 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2040); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2042 = 11'h7ea == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2041); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2043 = 11'h7eb == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2042); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2044 = 11'h7ec == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2043); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2045 = 11'h7ed == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2044); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2046 = 11'h7ee == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2045); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2047 = 11'h7ef == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2046); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2048 = 11'h7f0 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2047); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2049 = 11'h7f1 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2048); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2050 = 11'h7f2 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2049); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2051 = 11'h7f3 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2050); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2052 = 11'h7f4 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2051); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2053 = 11'h7f5 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2052); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2054 = 11'h7f6 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2053); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2055 = 11'h7f7 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2054); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2056 = 11'h7f8 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2055); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2057 = 11'h7f9 == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2056); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2058 = 11'h7fa == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2057); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2059 = 11'h7fb == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2058); // @[Reg.scala 17:{22,22}]
  wire [4:0] _GEN_2060 = 11'h7fc == data2In_0[10:0] ? $signed(5'shb) : $signed(_GEN_2059); // @[Reg.scala 17:{22,22}]
  wire [9:0] _data3In2_T_1 = 5'shb * $signed(data2Count_0); // @[logarithm.scala 56:81]
  reg [9:0] data3In2_0; // @[Reg.scala 16:16]
  wire [9:0] _GEN_2067 = {{5{data3In1_0[4]}},data3In1_0}; // @[logarithm.scala 58:71]
  wire [9:0] _data4_T_2 = $signed(_GEN_2067) + $signed(data3In2_0); // @[logarithm.scala 58:71]
  reg [9:0] data4_0; // @[Reg.scala 16:16]
  PipelineHsk_2 hsk ( // @[logarithm.scala 19:21]
    .clock(hsk_clock),
    .reset(hsk_reset),
    .io_validPre(hsk_io_validPre),
    .io_readyPre(hsk_io_readyPre),
    .io_lastPre(hsk_io_lastPre),
    .io_validNxt(hsk_io_validNxt),
    .io_readyNxt(hsk_io_readyNxt),
    .io_regen_0(hsk_io_regen_0),
    .io_regen_1(hsk_io_regen_1),
    .io_regen_2(hsk_io_regen_2),
    .io_regen_3(hsk_io_regen_3),
    .io_lastNxt(hsk_io_lastNxt)
  );
  assign io_output_valid = hsk_io_validNxt; // @[logarithm.scala 23:21]
  assign io_output_bits_x_0 = data4_0[7:0]; // @[logarithm.scala 59:22]
  assign hsk_clock = clock;
  assign hsk_reset = reset;
  assign hsk_io_validPre = io_input_valid; // @[logarithm.scala 20:21]
  assign hsk_io_lastPre = io_input_bits_last; // @[logarithm.scala 22:20]
  assign hsk_io_readyNxt = io_output_ready; // @[logarithm.scala 24:21]
  always @(posedge clock) begin
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_0 <= lod_0_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_1 <= lod_0_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_2 <= lod_0_2; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_3 <= lod_0_3; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_4 <= lod_0_4; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_5 <= lod_0_5; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_6 <= lod_0_6; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_7 <= lod_0_7; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_8 <= lod_0_8; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_9 <= lod_0_9; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_10 <= lod_0_10; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_11 <= lod_0_11; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1Lod_0_12 <= lod_0_12; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      data1In_0 <= io_input_bits_x_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2In_0 <= data2InMux_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_1) begin // @[Reg.scala 17:18]
      data2Count_0 <= data2CountMux_0; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_2) begin // @[Reg.scala 17:18]
      if (11'h7ff == data2In_0[10:0]) begin // @[Reg.scala 17:22]
        data3In1_0 <= 5'shb; // @[Reg.scala 17:22]
      end else if (11'h7fe == data2In_0[10:0]) begin // @[Reg.scala 17:22]
        data3In1_0 <= 5'shb; // @[Reg.scala 17:22]
      end else if (11'h7fd == data2In_0[10:0]) begin // @[Reg.scala 17:22]
        data3In1_0 <= 5'shb; // @[Reg.scala 17:22]
      end else begin
        data3In1_0 <= _GEN_2060;
      end
    end
    if (hsk_io_regen_2) begin // @[Reg.scala 17:18]
      data3In2_0 <= _data3In2_T_1; // @[Reg.scala 17:22]
    end
    if (hsk_io_regen_3) begin // @[Reg.scala 17:18]
      data4_0 <= _data4_T_2; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data1Lod_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  data1Lod_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data1Lod_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data1Lod_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  data1Lod_0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  data1Lod_0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  data1Lod_0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  data1Lod_0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  data1Lod_0_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  data1Lod_0_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  data1Lod_0_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  data1Lod_0_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  data1Lod_0_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  data1In_0 = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  data2In_0 = _RAND_14[11:0];
  _RAND_15 = {1{`RANDOM}};
  data2Count_0 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  data3In1_0 = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  data3In2_0 = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  data4_0 = _RAND_18[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Hsknto1(
  output       io_input_0_ready,
  input        io_input_0_valid,
  input  [7:0] io_input_0_bits_x_0,
  input  [7:0] io_input_0_bits_x_1,
  input  [7:0] io_input_0_bits_x_2,
  input  [7:0] io_input_0_bits_x_3,
  input  [7:0] io_input_0_bits_x_4,
  input  [7:0] io_input_0_bits_x_5,
  input  [7:0] io_input_0_bits_x_6,
  input  [7:0] io_input_0_bits_x_7,
  input  [7:0] io_input_0_bits_x_8,
  input  [7:0] io_input_0_bits_x_9,
  input  [7:0] io_input_0_bits_x_10,
  input  [7:0] io_input_0_bits_x_11,
  input  [7:0] io_input_0_bits_x_12,
  input  [7:0] io_input_0_bits_x_13,
  input  [7:0] io_input_0_bits_x_14,
  input  [7:0] io_input_0_bits_x_15,
  input        io_input_0_bits_last,
  output       io_input_1_ready,
  input        io_input_1_valid,
  input  [7:0] io_input_1_bits_x_0,
  input  [7:0] io_input_1_bits_x_1,
  input  [7:0] io_input_1_bits_x_2,
  input  [7:0] io_input_1_bits_x_3,
  input  [7:0] io_input_1_bits_x_4,
  input  [7:0] io_input_1_bits_x_5,
  input  [7:0] io_input_1_bits_x_6,
  input  [7:0] io_input_1_bits_x_7,
  input  [7:0] io_input_1_bits_x_8,
  input  [7:0] io_input_1_bits_x_9,
  input  [7:0] io_input_1_bits_x_10,
  input  [7:0] io_input_1_bits_x_11,
  input  [7:0] io_input_1_bits_x_12,
  input  [7:0] io_input_1_bits_x_13,
  input  [7:0] io_input_1_bits_x_14,
  input  [7:0] io_input_1_bits_x_15,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_0_x_0,
  output [7:0] io_output_bits_0_x_1,
  output [7:0] io_output_bits_0_x_2,
  output [7:0] io_output_bits_0_x_3,
  output [7:0] io_output_bits_0_x_4,
  output [7:0] io_output_bits_0_x_5,
  output [7:0] io_output_bits_0_x_6,
  output [7:0] io_output_bits_0_x_7,
  output [7:0] io_output_bits_0_x_8,
  output [7:0] io_output_bits_0_x_9,
  output [7:0] io_output_bits_0_x_10,
  output [7:0] io_output_bits_0_x_11,
  output [7:0] io_output_bits_0_x_12,
  output [7:0] io_output_bits_0_x_13,
  output [7:0] io_output_bits_0_x_14,
  output [7:0] io_output_bits_0_x_15,
  output       io_output_bits_0_last,
  output [7:0] io_output_bits_1_x_0,
  output [7:0] io_output_bits_1_x_1,
  output [7:0] io_output_bits_1_x_2,
  output [7:0] io_output_bits_1_x_3,
  output [7:0] io_output_bits_1_x_4,
  output [7:0] io_output_bits_1_x_5,
  output [7:0] io_output_bits_1_x_6,
  output [7:0] io_output_bits_1_x_7,
  output [7:0] io_output_bits_1_x_8,
  output [7:0] io_output_bits_1_x_9,
  output [7:0] io_output_bits_1_x_10,
  output [7:0] io_output_bits_1_x_11,
  output [7:0] io_output_bits_1_x_12,
  output [7:0] io_output_bits_1_x_13,
  output [7:0] io_output_bits_1_x_14,
  output [7:0] io_output_bits_1_x_15
);
  assign io_input_0_ready = io_output_ready & (~io_input_0_valid | io_input_1_valid); // @[hsknto1.scala 14:73]
  assign io_input_1_ready = io_output_ready & (~io_input_1_valid | io_input_0_valid); // @[hsknto1.scala 14:73]
  assign io_output_valid = io_input_0_valid & io_input_1_valid; // @[hsknto1.scala 12:58]
  assign io_output_bits_0_x_0 = io_input_0_bits_x_0; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_1 = io_input_0_bits_x_1; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_2 = io_input_0_bits_x_2; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_3 = io_input_0_bits_x_3; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_4 = io_input_0_bits_x_4; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_5 = io_input_0_bits_x_5; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_6 = io_input_0_bits_x_6; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_7 = io_input_0_bits_x_7; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_8 = io_input_0_bits_x_8; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_9 = io_input_0_bits_x_9; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_10 = io_input_0_bits_x_10; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_11 = io_input_0_bits_x_11; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_12 = io_input_0_bits_x_12; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_13 = io_input_0_bits_x_13; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_14 = io_input_0_bits_x_14; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_x_15 = io_input_0_bits_x_15; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_last = io_input_0_bits_last; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_0 = io_input_1_bits_x_0; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_1 = io_input_1_bits_x_1; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_2 = io_input_1_bits_x_2; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_3 = io_input_1_bits_x_3; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_4 = io_input_1_bits_x_4; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_5 = io_input_1_bits_x_5; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_6 = io_input_1_bits_x_6; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_7 = io_input_1_bits_x_7; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_8 = io_input_1_bits_x_8; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_9 = io_input_1_bits_x_9; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_10 = io_input_1_bits_x_10; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_11 = io_input_1_bits_x_11; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_12 = io_input_1_bits_x_12; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_13 = io_input_1_bits_x_13; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_14 = io_input_1_bits_x_14; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_15 = io_input_1_bits_x_15; // @[hsknto1.scala 13:55]
endmodule
module Softmax(
  input        clock,
  input        reset,
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_x_0,
  input  [7:0] io_input_bits_x_1,
  input  [7:0] io_input_bits_x_2,
  input  [7:0] io_input_bits_x_3,
  input  [7:0] io_input_bits_x_4,
  input  [7:0] io_input_bits_x_5,
  input  [7:0] io_input_bits_x_6,
  input  [7:0] io_input_bits_x_7,
  input  [7:0] io_input_bits_x_8,
  input  [7:0] io_input_bits_x_9,
  input  [7:0] io_input_bits_x_10,
  input  [7:0] io_input_bits_x_11,
  input  [7:0] io_input_bits_x_12,
  input  [7:0] io_input_bits_x_13,
  input  [7:0] io_input_bits_x_14,
  input  [7:0] io_input_bits_x_15,
  input        io_input_bits_last,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_x_0,
  output [7:0] io_output_bits_x_1,
  output [7:0] io_output_bits_x_2,
  output [7:0] io_output_bits_x_3,
  output [7:0] io_output_bits_x_4,
  output [7:0] io_output_bits_x_5,
  output [7:0] io_output_bits_x_6,
  output [7:0] io_output_bits_x_7,
  output [7:0] io_output_bits_x_8,
  output [7:0] io_output_bits_x_9,
  output [7:0] io_output_bits_x_10,
  output [7:0] io_output_bits_x_11,
  output [7:0] io_output_bits_x_12,
  output [7:0] io_output_bits_x_13,
  output [7:0] io_output_bits_x_14,
  output [7:0] io_output_bits_x_15,
  output       io_output_bits_last,
  input        rst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  exponentArray_clock; // @[softmax.scala 38:35]
  wire  exponentArray_reset; // @[softmax.scala 38:35]
  wire  exponentArray_io_input_ready; // @[softmax.scala 38:35]
  wire  exponentArray_io_input_valid; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_0; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_1; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_2; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_3; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_4; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_5; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_6; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_7; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_8; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_9; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_10; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_11; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_12; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_13; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_14; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_input_bits_x_15; // @[softmax.scala 38:35]
  wire  exponentArray_io_input_bits_last; // @[softmax.scala 38:35]
  wire  exponentArray_io_output_ready; // @[softmax.scala 38:35]
  wire  exponentArray_io_output_valid; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_0; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_1; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_2; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_3; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_4; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_5; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_6; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_7; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_8; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_9; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_10; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_11; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_12; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_13; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_14; // @[softmax.scala 38:35]
  wire [7:0] exponentArray_io_output_bits_x_15; // @[softmax.scala 38:35]
  wire  exponentArray_io_output_bits_last; // @[softmax.scala 38:35]
  wire  exponentArrayInHsk_io_input_ready; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_input_valid; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_0; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_1; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_2; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_3; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_4; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_5; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_6; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_7; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_8; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_9; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_10; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_11; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_12; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_13; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_14; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_0_x_15; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_input_bits_0_last; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_0; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_1; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_2; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_3; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_4; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_5; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_6; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_7; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_8; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_9; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_10; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_11; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_12; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_13; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_14; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_input_bits_1_x_15; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_input_bits_1_last; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_output_0_ready; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_output_0_valid; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_0; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_1; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_2; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_3; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_4; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_5; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_6; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_7; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_8; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_9; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_10; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_11; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_12; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_13; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_14; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_0_bits_x_15; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_output_0_bits_last; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_output_1_ready; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_output_1_valid; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_0; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_1; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_2; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_3; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_4; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_5; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_6; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_7; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_8; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_9; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_10; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_11; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_12; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_13; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_14; // @[softmax.scala 39:40]
  wire [7:0] exponentArrayInHsk_io_output_1_bits_x_15; // @[softmax.scala 39:40]
  wire  exponentArrayInHsk_io_output_1_bits_last; // @[softmax.scala 39:40]
  wire  exponentArrayInMux_io_input_0_ready; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_input_0_valid; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_0; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_1; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_2; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_3; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_4; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_5; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_6; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_7; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_8; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_9; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_10; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_11; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_12; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_13; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_14; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_0_bits_x_15; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_input_0_bits_last; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_input_1_ready; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_input_1_valid; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_0; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_1; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_2; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_3; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_4; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_5; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_6; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_7; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_8; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_9; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_10; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_11; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_12; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_13; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_14; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_input_1_bits_x_15; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_input_1_bits_last; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_sel; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_output_ready; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_output_valid; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_0; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_1; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_2; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_3; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_4; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_5; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_6; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_7; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_8; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_9; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_10; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_11; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_12; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_13; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_14; // @[softmax.scala 40:40]
  wire [7:0] exponentArrayInMux_io_output_bits_x_15; // @[softmax.scala 40:40]
  wire  exponentArrayInMux_io_output_bits_last; // @[softmax.scala 40:40]
  wire  exponentArrayOutMux_io_input_ready; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_input_valid; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_0; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_1; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_2; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_3; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_4; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_5; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_6; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_7; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_8; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_9; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_10; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_11; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_12; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_13; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_14; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_input_bits_x_15; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_input_bits_last; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_sel; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_output_0_ready; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_output_0_valid; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_0; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_1; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_2; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_3; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_4; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_5; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_6; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_7; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_8; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_9; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_10; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_11; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_12; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_13; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_14; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_0_bits_x_15; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_output_0_bits_last; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_output_1_ready; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_output_1_valid; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_0; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_1; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_2; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_3; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_4; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_5; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_6; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_7; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_8; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_9; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_10; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_11; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_12; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_13; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_14; // @[softmax.scala 41:41]
  wire [7:0] exponentArrayOutMux_io_output_1_bits_x_15; // @[softmax.scala 41:41]
  wire  exponentArrayOutMux_io_output_1_bits_last; // @[softmax.scala 41:41]
  wire  queue_clock; // @[softmax.scala 42:27]
  wire  queue_reset; // @[softmax.scala 42:27]
  wire  queue_io_enq_ready; // @[softmax.scala 42:27]
  wire  queue_io_enq_valid; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_0; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_1; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_2; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_3; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_4; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_5; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_6; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_7; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_8; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_9; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_10; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_11; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_12; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_13; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_14; // @[softmax.scala 42:27]
  wire [7:0] queue_io_enq_bits_x_15; // @[softmax.scala 42:27]
  wire  queue_io_enq_bits_last; // @[softmax.scala 42:27]
  wire  queue_io_deq_ready; // @[softmax.scala 42:27]
  wire  queue_io_deq_valid; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_0; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_1; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_2; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_3; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_4; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_5; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_6; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_7; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_8; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_9; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_10; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_11; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_12; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_13; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_14; // @[softmax.scala 42:27]
  wire [7:0] queue_io_deq_bits_x_15; // @[softmax.scala 42:27]
  wire  queue_io_deq_bits_last; // @[softmax.scala 42:27]
  wire  adder_clock; // @[softmax.scala 43:27]
  wire  adder_reset; // @[softmax.scala 43:27]
  wire  adder_io_input_ready; // @[softmax.scala 43:27]
  wire  adder_io_input_valid; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_0; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_1; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_2; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_3; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_4; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_5; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_6; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_7; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_8; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_9; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_10; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_11; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_12; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_13; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_14; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_15; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_16; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_17; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_18; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_19; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_20; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_21; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_22; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_23; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_24; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_25; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_26; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_27; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_28; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_29; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_30; // @[softmax.scala 43:27]
  wire [7:0] adder_io_input_bits_x_31; // @[softmax.scala 43:27]
  wire  adder_io_input_bits_last; // @[softmax.scala 43:27]
  wire  adder_io_output_ready; // @[softmax.scala 43:27]
  wire  adder_io_output_valid; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_0; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_1; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_2; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_3; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_4; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_5; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_6; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_7; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_8; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_9; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_10; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_11; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_12; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_13; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_14; // @[softmax.scala 43:27]
  wire [7:0] adder_io_output_bits_x_15; // @[softmax.scala 43:27]
  wire  adder_io_output_bits_last; // @[softmax.scala 43:27]
  wire  adderTree_clock; // @[softmax.scala 44:31]
  wire  adderTree_reset; // @[softmax.scala 44:31]
  wire  adderTree_io_input_ready; // @[softmax.scala 44:31]
  wire  adderTree_io_input_valid; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_0; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_1; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_2; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_3; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_4; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_5; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_6; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_7; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_8; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_9; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_10; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_11; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_12; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_13; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_14; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_input_bits_x_15; // @[softmax.scala 44:31]
  wire  adderTree_io_input_bits_last; // @[softmax.scala 44:31]
  wire  adderTree_io_output_valid; // @[softmax.scala 44:31]
  wire [11:0] adderTree_io_output_bits_x_0; // @[softmax.scala 44:31]
  wire  adderTree_io_output_bits_last; // @[softmax.scala 44:31]
  wire  accumulator_clock; // @[softmax.scala 45:33]
  wire  accumulator_reset; // @[softmax.scala 45:33]
  wire  accumulator_io_input_ready; // @[softmax.scala 45:33]
  wire  accumulator_io_input_valid; // @[softmax.scala 45:33]
  wire [11:0] accumulator_io_input_bits_x_0; // @[softmax.scala 45:33]
  wire  accumulator_io_input_bits_last; // @[softmax.scala 45:33]
  wire  accumulator_io_output_valid; // @[softmax.scala 45:33]
  wire [11:0] accumulator_io_output_bits_x_0; // @[softmax.scala 45:33]
  wire  accumulator_io_output_bits_last; // @[softmax.scala 45:33]
  wire  logarithm_clock; // @[softmax.scala 46:31]
  wire  logarithm_reset; // @[softmax.scala 46:31]
  wire  logarithm_io_input_valid; // @[softmax.scala 46:31]
  wire [11:0] logarithm_io_input_bits_x_0; // @[softmax.scala 46:31]
  wire  logarithm_io_input_bits_last; // @[softmax.scala 46:31]
  wire  logarithm_io_output_ready; // @[softmax.scala 46:31]
  wire  logarithm_io_output_valid; // @[softmax.scala 46:31]
  wire [7:0] logarithm_io_output_bits_x_0; // @[softmax.scala 46:31]
  wire  queueOutHsk_io_input_0_ready; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_input_0_valid; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_0; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_1; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_2; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_3; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_4; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_5; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_6; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_7; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_8; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_9; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_10; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_11; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_12; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_13; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_14; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_0_bits_x_15; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_input_0_bits_last; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_input_1_ready; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_input_1_valid; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_0; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_1; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_2; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_3; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_4; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_5; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_6; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_7; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_8; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_9; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_10; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_11; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_12; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_13; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_14; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_input_1_bits_x_15; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_output_ready; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_output_valid; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_0; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_1; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_2; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_3; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_4; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_5; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_6; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_7; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_8; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_9; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_10; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_11; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_12; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_13; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_14; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_0_x_15; // @[softmax.scala 47:33]
  wire  queueOutHsk_io_output_bits_0_last; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_0; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_1; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_2; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_3; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_4; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_5; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_6; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_7; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_8; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_9; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_10; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_11; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_12; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_13; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_14; // @[softmax.scala 47:33]
  wire [7:0] queueOutHsk_io_output_bits_1_x_15; // @[softmax.scala 47:33]
  reg  inPathSel; // @[Reg.scala 28:20]
  wire  inPathSelEn = exponentArray_io_input_valid & exponentArray_io_input_ready & exponentArray_io_input_bits_last; // @[softmax.scala 70:81]
  wire  inPathSelNxt = ~inPathSel; // @[softmax.scala 34:25]
  reg  outPathSel; // @[Reg.scala 28:20]
  wire  outPathSelEn = exponentArray_io_output_valid & exponentArray_io_output_ready & exponentArray_io_output_bits_last
    ; // @[softmax.scala 72:84]
  wire  outPathSelNxt = ~outPathSel; // @[softmax.scala 35:26]
  Exponent exponentArray ( // @[softmax.scala 38:35]
    .clock(exponentArray_clock),
    .reset(exponentArray_reset),
    .io_input_ready(exponentArray_io_input_ready),
    .io_input_valid(exponentArray_io_input_valid),
    .io_input_bits_x_0(exponentArray_io_input_bits_x_0),
    .io_input_bits_x_1(exponentArray_io_input_bits_x_1),
    .io_input_bits_x_2(exponentArray_io_input_bits_x_2),
    .io_input_bits_x_3(exponentArray_io_input_bits_x_3),
    .io_input_bits_x_4(exponentArray_io_input_bits_x_4),
    .io_input_bits_x_5(exponentArray_io_input_bits_x_5),
    .io_input_bits_x_6(exponentArray_io_input_bits_x_6),
    .io_input_bits_x_7(exponentArray_io_input_bits_x_7),
    .io_input_bits_x_8(exponentArray_io_input_bits_x_8),
    .io_input_bits_x_9(exponentArray_io_input_bits_x_9),
    .io_input_bits_x_10(exponentArray_io_input_bits_x_10),
    .io_input_bits_x_11(exponentArray_io_input_bits_x_11),
    .io_input_bits_x_12(exponentArray_io_input_bits_x_12),
    .io_input_bits_x_13(exponentArray_io_input_bits_x_13),
    .io_input_bits_x_14(exponentArray_io_input_bits_x_14),
    .io_input_bits_x_15(exponentArray_io_input_bits_x_15),
    .io_input_bits_last(exponentArray_io_input_bits_last),
    .io_output_ready(exponentArray_io_output_ready),
    .io_output_valid(exponentArray_io_output_valid),
    .io_output_bits_x_0(exponentArray_io_output_bits_x_0),
    .io_output_bits_x_1(exponentArray_io_output_bits_x_1),
    .io_output_bits_x_2(exponentArray_io_output_bits_x_2),
    .io_output_bits_x_3(exponentArray_io_output_bits_x_3),
    .io_output_bits_x_4(exponentArray_io_output_bits_x_4),
    .io_output_bits_x_5(exponentArray_io_output_bits_x_5),
    .io_output_bits_x_6(exponentArray_io_output_bits_x_6),
    .io_output_bits_x_7(exponentArray_io_output_bits_x_7),
    .io_output_bits_x_8(exponentArray_io_output_bits_x_8),
    .io_output_bits_x_9(exponentArray_io_output_bits_x_9),
    .io_output_bits_x_10(exponentArray_io_output_bits_x_10),
    .io_output_bits_x_11(exponentArray_io_output_bits_x_11),
    .io_output_bits_x_12(exponentArray_io_output_bits_x_12),
    .io_output_bits_x_13(exponentArray_io_output_bits_x_13),
    .io_output_bits_x_14(exponentArray_io_output_bits_x_14),
    .io_output_bits_x_15(exponentArray_io_output_bits_x_15),
    .io_output_bits_last(exponentArray_io_output_bits_last)
  );
  Hsk1ton exponentArrayInHsk ( // @[softmax.scala 39:40]
    .io_input_ready(exponentArrayInHsk_io_input_ready),
    .io_input_valid(exponentArrayInHsk_io_input_valid),
    .io_input_bits_0_x_0(exponentArrayInHsk_io_input_bits_0_x_0),
    .io_input_bits_0_x_1(exponentArrayInHsk_io_input_bits_0_x_1),
    .io_input_bits_0_x_2(exponentArrayInHsk_io_input_bits_0_x_2),
    .io_input_bits_0_x_3(exponentArrayInHsk_io_input_bits_0_x_3),
    .io_input_bits_0_x_4(exponentArrayInHsk_io_input_bits_0_x_4),
    .io_input_bits_0_x_5(exponentArrayInHsk_io_input_bits_0_x_5),
    .io_input_bits_0_x_6(exponentArrayInHsk_io_input_bits_0_x_6),
    .io_input_bits_0_x_7(exponentArrayInHsk_io_input_bits_0_x_7),
    .io_input_bits_0_x_8(exponentArrayInHsk_io_input_bits_0_x_8),
    .io_input_bits_0_x_9(exponentArrayInHsk_io_input_bits_0_x_9),
    .io_input_bits_0_x_10(exponentArrayInHsk_io_input_bits_0_x_10),
    .io_input_bits_0_x_11(exponentArrayInHsk_io_input_bits_0_x_11),
    .io_input_bits_0_x_12(exponentArrayInHsk_io_input_bits_0_x_12),
    .io_input_bits_0_x_13(exponentArrayInHsk_io_input_bits_0_x_13),
    .io_input_bits_0_x_14(exponentArrayInHsk_io_input_bits_0_x_14),
    .io_input_bits_0_x_15(exponentArrayInHsk_io_input_bits_0_x_15),
    .io_input_bits_0_last(exponentArrayInHsk_io_input_bits_0_last),
    .io_input_bits_1_x_0(exponentArrayInHsk_io_input_bits_1_x_0),
    .io_input_bits_1_x_1(exponentArrayInHsk_io_input_bits_1_x_1),
    .io_input_bits_1_x_2(exponentArrayInHsk_io_input_bits_1_x_2),
    .io_input_bits_1_x_3(exponentArrayInHsk_io_input_bits_1_x_3),
    .io_input_bits_1_x_4(exponentArrayInHsk_io_input_bits_1_x_4),
    .io_input_bits_1_x_5(exponentArrayInHsk_io_input_bits_1_x_5),
    .io_input_bits_1_x_6(exponentArrayInHsk_io_input_bits_1_x_6),
    .io_input_bits_1_x_7(exponentArrayInHsk_io_input_bits_1_x_7),
    .io_input_bits_1_x_8(exponentArrayInHsk_io_input_bits_1_x_8),
    .io_input_bits_1_x_9(exponentArrayInHsk_io_input_bits_1_x_9),
    .io_input_bits_1_x_10(exponentArrayInHsk_io_input_bits_1_x_10),
    .io_input_bits_1_x_11(exponentArrayInHsk_io_input_bits_1_x_11),
    .io_input_bits_1_x_12(exponentArrayInHsk_io_input_bits_1_x_12),
    .io_input_bits_1_x_13(exponentArrayInHsk_io_input_bits_1_x_13),
    .io_input_bits_1_x_14(exponentArrayInHsk_io_input_bits_1_x_14),
    .io_input_bits_1_x_15(exponentArrayInHsk_io_input_bits_1_x_15),
    .io_input_bits_1_last(exponentArrayInHsk_io_input_bits_1_last),
    .io_output_0_ready(exponentArrayInHsk_io_output_0_ready),
    .io_output_0_valid(exponentArrayInHsk_io_output_0_valid),
    .io_output_0_bits_x_0(exponentArrayInHsk_io_output_0_bits_x_0),
    .io_output_0_bits_x_1(exponentArrayInHsk_io_output_0_bits_x_1),
    .io_output_0_bits_x_2(exponentArrayInHsk_io_output_0_bits_x_2),
    .io_output_0_bits_x_3(exponentArrayInHsk_io_output_0_bits_x_3),
    .io_output_0_bits_x_4(exponentArrayInHsk_io_output_0_bits_x_4),
    .io_output_0_bits_x_5(exponentArrayInHsk_io_output_0_bits_x_5),
    .io_output_0_bits_x_6(exponentArrayInHsk_io_output_0_bits_x_6),
    .io_output_0_bits_x_7(exponentArrayInHsk_io_output_0_bits_x_7),
    .io_output_0_bits_x_8(exponentArrayInHsk_io_output_0_bits_x_8),
    .io_output_0_bits_x_9(exponentArrayInHsk_io_output_0_bits_x_9),
    .io_output_0_bits_x_10(exponentArrayInHsk_io_output_0_bits_x_10),
    .io_output_0_bits_x_11(exponentArrayInHsk_io_output_0_bits_x_11),
    .io_output_0_bits_x_12(exponentArrayInHsk_io_output_0_bits_x_12),
    .io_output_0_bits_x_13(exponentArrayInHsk_io_output_0_bits_x_13),
    .io_output_0_bits_x_14(exponentArrayInHsk_io_output_0_bits_x_14),
    .io_output_0_bits_x_15(exponentArrayInHsk_io_output_0_bits_x_15),
    .io_output_0_bits_last(exponentArrayInHsk_io_output_0_bits_last),
    .io_output_1_ready(exponentArrayInHsk_io_output_1_ready),
    .io_output_1_valid(exponentArrayInHsk_io_output_1_valid),
    .io_output_1_bits_x_0(exponentArrayInHsk_io_output_1_bits_x_0),
    .io_output_1_bits_x_1(exponentArrayInHsk_io_output_1_bits_x_1),
    .io_output_1_bits_x_2(exponentArrayInHsk_io_output_1_bits_x_2),
    .io_output_1_bits_x_3(exponentArrayInHsk_io_output_1_bits_x_3),
    .io_output_1_bits_x_4(exponentArrayInHsk_io_output_1_bits_x_4),
    .io_output_1_bits_x_5(exponentArrayInHsk_io_output_1_bits_x_5),
    .io_output_1_bits_x_6(exponentArrayInHsk_io_output_1_bits_x_6),
    .io_output_1_bits_x_7(exponentArrayInHsk_io_output_1_bits_x_7),
    .io_output_1_bits_x_8(exponentArrayInHsk_io_output_1_bits_x_8),
    .io_output_1_bits_x_9(exponentArrayInHsk_io_output_1_bits_x_9),
    .io_output_1_bits_x_10(exponentArrayInHsk_io_output_1_bits_x_10),
    .io_output_1_bits_x_11(exponentArrayInHsk_io_output_1_bits_x_11),
    .io_output_1_bits_x_12(exponentArrayInHsk_io_output_1_bits_x_12),
    .io_output_1_bits_x_13(exponentArrayInHsk_io_output_1_bits_x_13),
    .io_output_1_bits_x_14(exponentArrayInHsk_io_output_1_bits_x_14),
    .io_output_1_bits_x_15(exponentArrayInHsk_io_output_1_bits_x_15),
    .io_output_1_bits_last(exponentArrayInHsk_io_output_1_bits_last)
  );
  Arbiternto1 exponentArrayInMux ( // @[softmax.scala 40:40]
    .io_input_0_ready(exponentArrayInMux_io_input_0_ready),
    .io_input_0_valid(exponentArrayInMux_io_input_0_valid),
    .io_input_0_bits_x_0(exponentArrayInMux_io_input_0_bits_x_0),
    .io_input_0_bits_x_1(exponentArrayInMux_io_input_0_bits_x_1),
    .io_input_0_bits_x_2(exponentArrayInMux_io_input_0_bits_x_2),
    .io_input_0_bits_x_3(exponentArrayInMux_io_input_0_bits_x_3),
    .io_input_0_bits_x_4(exponentArrayInMux_io_input_0_bits_x_4),
    .io_input_0_bits_x_5(exponentArrayInMux_io_input_0_bits_x_5),
    .io_input_0_bits_x_6(exponentArrayInMux_io_input_0_bits_x_6),
    .io_input_0_bits_x_7(exponentArrayInMux_io_input_0_bits_x_7),
    .io_input_0_bits_x_8(exponentArrayInMux_io_input_0_bits_x_8),
    .io_input_0_bits_x_9(exponentArrayInMux_io_input_0_bits_x_9),
    .io_input_0_bits_x_10(exponentArrayInMux_io_input_0_bits_x_10),
    .io_input_0_bits_x_11(exponentArrayInMux_io_input_0_bits_x_11),
    .io_input_0_bits_x_12(exponentArrayInMux_io_input_0_bits_x_12),
    .io_input_0_bits_x_13(exponentArrayInMux_io_input_0_bits_x_13),
    .io_input_0_bits_x_14(exponentArrayInMux_io_input_0_bits_x_14),
    .io_input_0_bits_x_15(exponentArrayInMux_io_input_0_bits_x_15),
    .io_input_0_bits_last(exponentArrayInMux_io_input_0_bits_last),
    .io_input_1_ready(exponentArrayInMux_io_input_1_ready),
    .io_input_1_valid(exponentArrayInMux_io_input_1_valid),
    .io_input_1_bits_x_0(exponentArrayInMux_io_input_1_bits_x_0),
    .io_input_1_bits_x_1(exponentArrayInMux_io_input_1_bits_x_1),
    .io_input_1_bits_x_2(exponentArrayInMux_io_input_1_bits_x_2),
    .io_input_1_bits_x_3(exponentArrayInMux_io_input_1_bits_x_3),
    .io_input_1_bits_x_4(exponentArrayInMux_io_input_1_bits_x_4),
    .io_input_1_bits_x_5(exponentArrayInMux_io_input_1_bits_x_5),
    .io_input_1_bits_x_6(exponentArrayInMux_io_input_1_bits_x_6),
    .io_input_1_bits_x_7(exponentArrayInMux_io_input_1_bits_x_7),
    .io_input_1_bits_x_8(exponentArrayInMux_io_input_1_bits_x_8),
    .io_input_1_bits_x_9(exponentArrayInMux_io_input_1_bits_x_9),
    .io_input_1_bits_x_10(exponentArrayInMux_io_input_1_bits_x_10),
    .io_input_1_bits_x_11(exponentArrayInMux_io_input_1_bits_x_11),
    .io_input_1_bits_x_12(exponentArrayInMux_io_input_1_bits_x_12),
    .io_input_1_bits_x_13(exponentArrayInMux_io_input_1_bits_x_13),
    .io_input_1_bits_x_14(exponentArrayInMux_io_input_1_bits_x_14),
    .io_input_1_bits_x_15(exponentArrayInMux_io_input_1_bits_x_15),
    .io_input_1_bits_last(exponentArrayInMux_io_input_1_bits_last),
    .io_sel(exponentArrayInMux_io_sel),
    .io_output_ready(exponentArrayInMux_io_output_ready),
    .io_output_valid(exponentArrayInMux_io_output_valid),
    .io_output_bits_x_0(exponentArrayInMux_io_output_bits_x_0),
    .io_output_bits_x_1(exponentArrayInMux_io_output_bits_x_1),
    .io_output_bits_x_2(exponentArrayInMux_io_output_bits_x_2),
    .io_output_bits_x_3(exponentArrayInMux_io_output_bits_x_3),
    .io_output_bits_x_4(exponentArrayInMux_io_output_bits_x_4),
    .io_output_bits_x_5(exponentArrayInMux_io_output_bits_x_5),
    .io_output_bits_x_6(exponentArrayInMux_io_output_bits_x_6),
    .io_output_bits_x_7(exponentArrayInMux_io_output_bits_x_7),
    .io_output_bits_x_8(exponentArrayInMux_io_output_bits_x_8),
    .io_output_bits_x_9(exponentArrayInMux_io_output_bits_x_9),
    .io_output_bits_x_10(exponentArrayInMux_io_output_bits_x_10),
    .io_output_bits_x_11(exponentArrayInMux_io_output_bits_x_11),
    .io_output_bits_x_12(exponentArrayInMux_io_output_bits_x_12),
    .io_output_bits_x_13(exponentArrayInMux_io_output_bits_x_13),
    .io_output_bits_x_14(exponentArrayInMux_io_output_bits_x_14),
    .io_output_bits_x_15(exponentArrayInMux_io_output_bits_x_15),
    .io_output_bits_last(exponentArrayInMux_io_output_bits_last)
  );
  Arbiter1ton exponentArrayOutMux ( // @[softmax.scala 41:41]
    .io_input_ready(exponentArrayOutMux_io_input_ready),
    .io_input_valid(exponentArrayOutMux_io_input_valid),
    .io_input_bits_x_0(exponentArrayOutMux_io_input_bits_x_0),
    .io_input_bits_x_1(exponentArrayOutMux_io_input_bits_x_1),
    .io_input_bits_x_2(exponentArrayOutMux_io_input_bits_x_2),
    .io_input_bits_x_3(exponentArrayOutMux_io_input_bits_x_3),
    .io_input_bits_x_4(exponentArrayOutMux_io_input_bits_x_4),
    .io_input_bits_x_5(exponentArrayOutMux_io_input_bits_x_5),
    .io_input_bits_x_6(exponentArrayOutMux_io_input_bits_x_6),
    .io_input_bits_x_7(exponentArrayOutMux_io_input_bits_x_7),
    .io_input_bits_x_8(exponentArrayOutMux_io_input_bits_x_8),
    .io_input_bits_x_9(exponentArrayOutMux_io_input_bits_x_9),
    .io_input_bits_x_10(exponentArrayOutMux_io_input_bits_x_10),
    .io_input_bits_x_11(exponentArrayOutMux_io_input_bits_x_11),
    .io_input_bits_x_12(exponentArrayOutMux_io_input_bits_x_12),
    .io_input_bits_x_13(exponentArrayOutMux_io_input_bits_x_13),
    .io_input_bits_x_14(exponentArrayOutMux_io_input_bits_x_14),
    .io_input_bits_x_15(exponentArrayOutMux_io_input_bits_x_15),
    .io_input_bits_last(exponentArrayOutMux_io_input_bits_last),
    .io_sel(exponentArrayOutMux_io_sel),
    .io_output_0_ready(exponentArrayOutMux_io_output_0_ready),
    .io_output_0_valid(exponentArrayOutMux_io_output_0_valid),
    .io_output_0_bits_x_0(exponentArrayOutMux_io_output_0_bits_x_0),
    .io_output_0_bits_x_1(exponentArrayOutMux_io_output_0_bits_x_1),
    .io_output_0_bits_x_2(exponentArrayOutMux_io_output_0_bits_x_2),
    .io_output_0_bits_x_3(exponentArrayOutMux_io_output_0_bits_x_3),
    .io_output_0_bits_x_4(exponentArrayOutMux_io_output_0_bits_x_4),
    .io_output_0_bits_x_5(exponentArrayOutMux_io_output_0_bits_x_5),
    .io_output_0_bits_x_6(exponentArrayOutMux_io_output_0_bits_x_6),
    .io_output_0_bits_x_7(exponentArrayOutMux_io_output_0_bits_x_7),
    .io_output_0_bits_x_8(exponentArrayOutMux_io_output_0_bits_x_8),
    .io_output_0_bits_x_9(exponentArrayOutMux_io_output_0_bits_x_9),
    .io_output_0_bits_x_10(exponentArrayOutMux_io_output_0_bits_x_10),
    .io_output_0_bits_x_11(exponentArrayOutMux_io_output_0_bits_x_11),
    .io_output_0_bits_x_12(exponentArrayOutMux_io_output_0_bits_x_12),
    .io_output_0_bits_x_13(exponentArrayOutMux_io_output_0_bits_x_13),
    .io_output_0_bits_x_14(exponentArrayOutMux_io_output_0_bits_x_14),
    .io_output_0_bits_x_15(exponentArrayOutMux_io_output_0_bits_x_15),
    .io_output_0_bits_last(exponentArrayOutMux_io_output_0_bits_last),
    .io_output_1_ready(exponentArrayOutMux_io_output_1_ready),
    .io_output_1_valid(exponentArrayOutMux_io_output_1_valid),
    .io_output_1_bits_x_0(exponentArrayOutMux_io_output_1_bits_x_0),
    .io_output_1_bits_x_1(exponentArrayOutMux_io_output_1_bits_x_1),
    .io_output_1_bits_x_2(exponentArrayOutMux_io_output_1_bits_x_2),
    .io_output_1_bits_x_3(exponentArrayOutMux_io_output_1_bits_x_3),
    .io_output_1_bits_x_4(exponentArrayOutMux_io_output_1_bits_x_4),
    .io_output_1_bits_x_5(exponentArrayOutMux_io_output_1_bits_x_5),
    .io_output_1_bits_x_6(exponentArrayOutMux_io_output_1_bits_x_6),
    .io_output_1_bits_x_7(exponentArrayOutMux_io_output_1_bits_x_7),
    .io_output_1_bits_x_8(exponentArrayOutMux_io_output_1_bits_x_8),
    .io_output_1_bits_x_9(exponentArrayOutMux_io_output_1_bits_x_9),
    .io_output_1_bits_x_10(exponentArrayOutMux_io_output_1_bits_x_10),
    .io_output_1_bits_x_11(exponentArrayOutMux_io_output_1_bits_x_11),
    .io_output_1_bits_x_12(exponentArrayOutMux_io_output_1_bits_x_12),
    .io_output_1_bits_x_13(exponentArrayOutMux_io_output_1_bits_x_13),
    .io_output_1_bits_x_14(exponentArrayOutMux_io_output_1_bits_x_14),
    .io_output_1_bits_x_15(exponentArrayOutMux_io_output_1_bits_x_15),
    .io_output_1_bits_last(exponentArrayOutMux_io_output_1_bits_last)
  );
  Queue queue ( // @[softmax.scala 42:27]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_x_0(queue_io_enq_bits_x_0),
    .io_enq_bits_x_1(queue_io_enq_bits_x_1),
    .io_enq_bits_x_2(queue_io_enq_bits_x_2),
    .io_enq_bits_x_3(queue_io_enq_bits_x_3),
    .io_enq_bits_x_4(queue_io_enq_bits_x_4),
    .io_enq_bits_x_5(queue_io_enq_bits_x_5),
    .io_enq_bits_x_6(queue_io_enq_bits_x_6),
    .io_enq_bits_x_7(queue_io_enq_bits_x_7),
    .io_enq_bits_x_8(queue_io_enq_bits_x_8),
    .io_enq_bits_x_9(queue_io_enq_bits_x_9),
    .io_enq_bits_x_10(queue_io_enq_bits_x_10),
    .io_enq_bits_x_11(queue_io_enq_bits_x_11),
    .io_enq_bits_x_12(queue_io_enq_bits_x_12),
    .io_enq_bits_x_13(queue_io_enq_bits_x_13),
    .io_enq_bits_x_14(queue_io_enq_bits_x_14),
    .io_enq_bits_x_15(queue_io_enq_bits_x_15),
    .io_enq_bits_last(queue_io_enq_bits_last),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_x_0(queue_io_deq_bits_x_0),
    .io_deq_bits_x_1(queue_io_deq_bits_x_1),
    .io_deq_bits_x_2(queue_io_deq_bits_x_2),
    .io_deq_bits_x_3(queue_io_deq_bits_x_3),
    .io_deq_bits_x_4(queue_io_deq_bits_x_4),
    .io_deq_bits_x_5(queue_io_deq_bits_x_5),
    .io_deq_bits_x_6(queue_io_deq_bits_x_6),
    .io_deq_bits_x_7(queue_io_deq_bits_x_7),
    .io_deq_bits_x_8(queue_io_deq_bits_x_8),
    .io_deq_bits_x_9(queue_io_deq_bits_x_9),
    .io_deq_bits_x_10(queue_io_deq_bits_x_10),
    .io_deq_bits_x_11(queue_io_deq_bits_x_11),
    .io_deq_bits_x_12(queue_io_deq_bits_x_12),
    .io_deq_bits_x_13(queue_io_deq_bits_x_13),
    .io_deq_bits_x_14(queue_io_deq_bits_x_14),
    .io_deq_bits_x_15(queue_io_deq_bits_x_15),
    .io_deq_bits_last(queue_io_deq_bits_last)
  );
  Adder2to1 adder ( // @[softmax.scala 43:27]
    .clock(adder_clock),
    .reset(adder_reset),
    .io_input_ready(adder_io_input_ready),
    .io_input_valid(adder_io_input_valid),
    .io_input_bits_x_0(adder_io_input_bits_x_0),
    .io_input_bits_x_1(adder_io_input_bits_x_1),
    .io_input_bits_x_2(adder_io_input_bits_x_2),
    .io_input_bits_x_3(adder_io_input_bits_x_3),
    .io_input_bits_x_4(adder_io_input_bits_x_4),
    .io_input_bits_x_5(adder_io_input_bits_x_5),
    .io_input_bits_x_6(adder_io_input_bits_x_6),
    .io_input_bits_x_7(adder_io_input_bits_x_7),
    .io_input_bits_x_8(adder_io_input_bits_x_8),
    .io_input_bits_x_9(adder_io_input_bits_x_9),
    .io_input_bits_x_10(adder_io_input_bits_x_10),
    .io_input_bits_x_11(adder_io_input_bits_x_11),
    .io_input_bits_x_12(adder_io_input_bits_x_12),
    .io_input_bits_x_13(adder_io_input_bits_x_13),
    .io_input_bits_x_14(adder_io_input_bits_x_14),
    .io_input_bits_x_15(adder_io_input_bits_x_15),
    .io_input_bits_x_16(adder_io_input_bits_x_16),
    .io_input_bits_x_17(adder_io_input_bits_x_17),
    .io_input_bits_x_18(adder_io_input_bits_x_18),
    .io_input_bits_x_19(adder_io_input_bits_x_19),
    .io_input_bits_x_20(adder_io_input_bits_x_20),
    .io_input_bits_x_21(adder_io_input_bits_x_21),
    .io_input_bits_x_22(adder_io_input_bits_x_22),
    .io_input_bits_x_23(adder_io_input_bits_x_23),
    .io_input_bits_x_24(adder_io_input_bits_x_24),
    .io_input_bits_x_25(adder_io_input_bits_x_25),
    .io_input_bits_x_26(adder_io_input_bits_x_26),
    .io_input_bits_x_27(adder_io_input_bits_x_27),
    .io_input_bits_x_28(adder_io_input_bits_x_28),
    .io_input_bits_x_29(adder_io_input_bits_x_29),
    .io_input_bits_x_30(adder_io_input_bits_x_30),
    .io_input_bits_x_31(adder_io_input_bits_x_31),
    .io_input_bits_last(adder_io_input_bits_last),
    .io_output_ready(adder_io_output_ready),
    .io_output_valid(adder_io_output_valid),
    .io_output_bits_x_0(adder_io_output_bits_x_0),
    .io_output_bits_x_1(adder_io_output_bits_x_1),
    .io_output_bits_x_2(adder_io_output_bits_x_2),
    .io_output_bits_x_3(adder_io_output_bits_x_3),
    .io_output_bits_x_4(adder_io_output_bits_x_4),
    .io_output_bits_x_5(adder_io_output_bits_x_5),
    .io_output_bits_x_6(adder_io_output_bits_x_6),
    .io_output_bits_x_7(adder_io_output_bits_x_7),
    .io_output_bits_x_8(adder_io_output_bits_x_8),
    .io_output_bits_x_9(adder_io_output_bits_x_9),
    .io_output_bits_x_10(adder_io_output_bits_x_10),
    .io_output_bits_x_11(adder_io_output_bits_x_11),
    .io_output_bits_x_12(adder_io_output_bits_x_12),
    .io_output_bits_x_13(adder_io_output_bits_x_13),
    .io_output_bits_x_14(adder_io_output_bits_x_14),
    .io_output_bits_x_15(adder_io_output_bits_x_15),
    .io_output_bits_last(adder_io_output_bits_last)
  );
  AdderTree adderTree ( // @[softmax.scala 44:31]
    .clock(adderTree_clock),
    .reset(adderTree_reset),
    .io_input_ready(adderTree_io_input_ready),
    .io_input_valid(adderTree_io_input_valid),
    .io_input_bits_x_0(adderTree_io_input_bits_x_0),
    .io_input_bits_x_1(adderTree_io_input_bits_x_1),
    .io_input_bits_x_2(adderTree_io_input_bits_x_2),
    .io_input_bits_x_3(adderTree_io_input_bits_x_3),
    .io_input_bits_x_4(adderTree_io_input_bits_x_4),
    .io_input_bits_x_5(adderTree_io_input_bits_x_5),
    .io_input_bits_x_6(adderTree_io_input_bits_x_6),
    .io_input_bits_x_7(adderTree_io_input_bits_x_7),
    .io_input_bits_x_8(adderTree_io_input_bits_x_8),
    .io_input_bits_x_9(adderTree_io_input_bits_x_9),
    .io_input_bits_x_10(adderTree_io_input_bits_x_10),
    .io_input_bits_x_11(adderTree_io_input_bits_x_11),
    .io_input_bits_x_12(adderTree_io_input_bits_x_12),
    .io_input_bits_x_13(adderTree_io_input_bits_x_13),
    .io_input_bits_x_14(adderTree_io_input_bits_x_14),
    .io_input_bits_x_15(adderTree_io_input_bits_x_15),
    .io_input_bits_last(adderTree_io_input_bits_last),
    .io_output_valid(adderTree_io_output_valid),
    .io_output_bits_x_0(adderTree_io_output_bits_x_0),
    .io_output_bits_last(adderTree_io_output_bits_last)
  );
  Accumulator2to1 accumulator ( // @[softmax.scala 45:33]
    .clock(accumulator_clock),
    .reset(accumulator_reset),
    .io_input_ready(accumulator_io_input_ready),
    .io_input_valid(accumulator_io_input_valid),
    .io_input_bits_x_0(accumulator_io_input_bits_x_0),
    .io_input_bits_last(accumulator_io_input_bits_last),
    .io_output_valid(accumulator_io_output_valid),
    .io_output_bits_x_0(accumulator_io_output_bits_x_0),
    .io_output_bits_last(accumulator_io_output_bits_last)
  );
  Logarithm logarithm ( // @[softmax.scala 46:31]
    .clock(logarithm_clock),
    .reset(logarithm_reset),
    .io_input_valid(logarithm_io_input_valid),
    .io_input_bits_x_0(logarithm_io_input_bits_x_0),
    .io_input_bits_last(logarithm_io_input_bits_last),
    .io_output_ready(logarithm_io_output_ready),
    .io_output_valid(logarithm_io_output_valid),
    .io_output_bits_x_0(logarithm_io_output_bits_x_0)
  );
  Hsknto1 queueOutHsk ( // @[softmax.scala 47:33]
    .io_input_0_ready(queueOutHsk_io_input_0_ready),
    .io_input_0_valid(queueOutHsk_io_input_0_valid),
    .io_input_0_bits_x_0(queueOutHsk_io_input_0_bits_x_0),
    .io_input_0_bits_x_1(queueOutHsk_io_input_0_bits_x_1),
    .io_input_0_bits_x_2(queueOutHsk_io_input_0_bits_x_2),
    .io_input_0_bits_x_3(queueOutHsk_io_input_0_bits_x_3),
    .io_input_0_bits_x_4(queueOutHsk_io_input_0_bits_x_4),
    .io_input_0_bits_x_5(queueOutHsk_io_input_0_bits_x_5),
    .io_input_0_bits_x_6(queueOutHsk_io_input_0_bits_x_6),
    .io_input_0_bits_x_7(queueOutHsk_io_input_0_bits_x_7),
    .io_input_0_bits_x_8(queueOutHsk_io_input_0_bits_x_8),
    .io_input_0_bits_x_9(queueOutHsk_io_input_0_bits_x_9),
    .io_input_0_bits_x_10(queueOutHsk_io_input_0_bits_x_10),
    .io_input_0_bits_x_11(queueOutHsk_io_input_0_bits_x_11),
    .io_input_0_bits_x_12(queueOutHsk_io_input_0_bits_x_12),
    .io_input_0_bits_x_13(queueOutHsk_io_input_0_bits_x_13),
    .io_input_0_bits_x_14(queueOutHsk_io_input_0_bits_x_14),
    .io_input_0_bits_x_15(queueOutHsk_io_input_0_bits_x_15),
    .io_input_0_bits_last(queueOutHsk_io_input_0_bits_last),
    .io_input_1_ready(queueOutHsk_io_input_1_ready),
    .io_input_1_valid(queueOutHsk_io_input_1_valid),
    .io_input_1_bits_x_0(queueOutHsk_io_input_1_bits_x_0),
    .io_input_1_bits_x_1(queueOutHsk_io_input_1_bits_x_1),
    .io_input_1_bits_x_2(queueOutHsk_io_input_1_bits_x_2),
    .io_input_1_bits_x_3(queueOutHsk_io_input_1_bits_x_3),
    .io_input_1_bits_x_4(queueOutHsk_io_input_1_bits_x_4),
    .io_input_1_bits_x_5(queueOutHsk_io_input_1_bits_x_5),
    .io_input_1_bits_x_6(queueOutHsk_io_input_1_bits_x_6),
    .io_input_1_bits_x_7(queueOutHsk_io_input_1_bits_x_7),
    .io_input_1_bits_x_8(queueOutHsk_io_input_1_bits_x_8),
    .io_input_1_bits_x_9(queueOutHsk_io_input_1_bits_x_9),
    .io_input_1_bits_x_10(queueOutHsk_io_input_1_bits_x_10),
    .io_input_1_bits_x_11(queueOutHsk_io_input_1_bits_x_11),
    .io_input_1_bits_x_12(queueOutHsk_io_input_1_bits_x_12),
    .io_input_1_bits_x_13(queueOutHsk_io_input_1_bits_x_13),
    .io_input_1_bits_x_14(queueOutHsk_io_input_1_bits_x_14),
    .io_input_1_bits_x_15(queueOutHsk_io_input_1_bits_x_15),
    .io_output_ready(queueOutHsk_io_output_ready),
    .io_output_valid(queueOutHsk_io_output_valid),
    .io_output_bits_0_x_0(queueOutHsk_io_output_bits_0_x_0),
    .io_output_bits_0_x_1(queueOutHsk_io_output_bits_0_x_1),
    .io_output_bits_0_x_2(queueOutHsk_io_output_bits_0_x_2),
    .io_output_bits_0_x_3(queueOutHsk_io_output_bits_0_x_3),
    .io_output_bits_0_x_4(queueOutHsk_io_output_bits_0_x_4),
    .io_output_bits_0_x_5(queueOutHsk_io_output_bits_0_x_5),
    .io_output_bits_0_x_6(queueOutHsk_io_output_bits_0_x_6),
    .io_output_bits_0_x_7(queueOutHsk_io_output_bits_0_x_7),
    .io_output_bits_0_x_8(queueOutHsk_io_output_bits_0_x_8),
    .io_output_bits_0_x_9(queueOutHsk_io_output_bits_0_x_9),
    .io_output_bits_0_x_10(queueOutHsk_io_output_bits_0_x_10),
    .io_output_bits_0_x_11(queueOutHsk_io_output_bits_0_x_11),
    .io_output_bits_0_x_12(queueOutHsk_io_output_bits_0_x_12),
    .io_output_bits_0_x_13(queueOutHsk_io_output_bits_0_x_13),
    .io_output_bits_0_x_14(queueOutHsk_io_output_bits_0_x_14),
    .io_output_bits_0_x_15(queueOutHsk_io_output_bits_0_x_15),
    .io_output_bits_0_last(queueOutHsk_io_output_bits_0_last),
    .io_output_bits_1_x_0(queueOutHsk_io_output_bits_1_x_0),
    .io_output_bits_1_x_1(queueOutHsk_io_output_bits_1_x_1),
    .io_output_bits_1_x_2(queueOutHsk_io_output_bits_1_x_2),
    .io_output_bits_1_x_3(queueOutHsk_io_output_bits_1_x_3),
    .io_output_bits_1_x_4(queueOutHsk_io_output_bits_1_x_4),
    .io_output_bits_1_x_5(queueOutHsk_io_output_bits_1_x_5),
    .io_output_bits_1_x_6(queueOutHsk_io_output_bits_1_x_6),
    .io_output_bits_1_x_7(queueOutHsk_io_output_bits_1_x_7),
    .io_output_bits_1_x_8(queueOutHsk_io_output_bits_1_x_8),
    .io_output_bits_1_x_9(queueOutHsk_io_output_bits_1_x_9),
    .io_output_bits_1_x_10(queueOutHsk_io_output_bits_1_x_10),
    .io_output_bits_1_x_11(queueOutHsk_io_output_bits_1_x_11),
    .io_output_bits_1_x_12(queueOutHsk_io_output_bits_1_x_12),
    .io_output_bits_1_x_13(queueOutHsk_io_output_bits_1_x_13),
    .io_output_bits_1_x_14(queueOutHsk_io_output_bits_1_x_14),
    .io_output_bits_1_x_15(queueOutHsk_io_output_bits_1_x_15)
  );
  assign io_input_ready = exponentArrayInHsk_io_input_ready; // @[port.scala 68:19]
  assign io_output_valid = exponentArrayOutMux_io_output_1_valid; // @[softmax.scala 59:42]
  assign io_output_bits_x_0 = exponentArrayOutMux_io_output_1_bits_x_0; // @[softmax.scala 59:42]
  assign io_output_bits_x_1 = exponentArrayOutMux_io_output_1_bits_x_1; // @[softmax.scala 59:42]
  assign io_output_bits_x_2 = exponentArrayOutMux_io_output_1_bits_x_2; // @[softmax.scala 59:42]
  assign io_output_bits_x_3 = exponentArrayOutMux_io_output_1_bits_x_3; // @[softmax.scala 59:42]
  assign io_output_bits_x_4 = exponentArrayOutMux_io_output_1_bits_x_4; // @[softmax.scala 59:42]
  assign io_output_bits_x_5 = exponentArrayOutMux_io_output_1_bits_x_5; // @[softmax.scala 59:42]
  assign io_output_bits_x_6 = exponentArrayOutMux_io_output_1_bits_x_6; // @[softmax.scala 59:42]
  assign io_output_bits_x_7 = exponentArrayOutMux_io_output_1_bits_x_7; // @[softmax.scala 59:42]
  assign io_output_bits_x_8 = exponentArrayOutMux_io_output_1_bits_x_8; // @[softmax.scala 59:42]
  assign io_output_bits_x_9 = exponentArrayOutMux_io_output_1_bits_x_9; // @[softmax.scala 59:42]
  assign io_output_bits_x_10 = exponentArrayOutMux_io_output_1_bits_x_10; // @[softmax.scala 59:42]
  assign io_output_bits_x_11 = exponentArrayOutMux_io_output_1_bits_x_11; // @[softmax.scala 59:42]
  assign io_output_bits_x_12 = exponentArrayOutMux_io_output_1_bits_x_12; // @[softmax.scala 59:42]
  assign io_output_bits_x_13 = exponentArrayOutMux_io_output_1_bits_x_13; // @[softmax.scala 59:42]
  assign io_output_bits_x_14 = exponentArrayOutMux_io_output_1_bits_x_14; // @[softmax.scala 59:42]
  assign io_output_bits_x_15 = exponentArrayOutMux_io_output_1_bits_x_15; // @[softmax.scala 59:42]
  assign io_output_bits_last = exponentArrayOutMux_io_output_1_bits_last; // @[softmax.scala 59:42]
  assign exponentArray_clock = clock;
  assign exponentArray_reset = rst;
  assign exponentArray_io_input_valid = exponentArrayInMux_io_output_valid; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_0 = exponentArrayInMux_io_output_bits_x_0; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_1 = exponentArrayInMux_io_output_bits_x_1; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_2 = exponentArrayInMux_io_output_bits_x_2; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_3 = exponentArrayInMux_io_output_bits_x_3; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_4 = exponentArrayInMux_io_output_bits_x_4; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_5 = exponentArrayInMux_io_output_bits_x_5; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_6 = exponentArrayInMux_io_output_bits_x_6; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_7 = exponentArrayInMux_io_output_bits_x_7; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_8 = exponentArrayInMux_io_output_bits_x_8; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_9 = exponentArrayInMux_io_output_bits_x_9; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_10 = exponentArrayInMux_io_output_bits_x_10; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_11 = exponentArrayInMux_io_output_bits_x_11; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_12 = exponentArrayInMux_io_output_bits_x_12; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_13 = exponentArrayInMux_io_output_bits_x_13; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_14 = exponentArrayInMux_io_output_bits_x_14; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_x_15 = exponentArrayInMux_io_output_bits_x_15; // @[softmax.scala 54:38]
  assign exponentArray_io_input_bits_last = exponentArrayInMux_io_output_bits_last; // @[softmax.scala 54:38]
  assign exponentArray_io_output_ready = exponentArrayOutMux_io_input_ready; // @[softmax.scala 57:33]
  assign exponentArrayInHsk_io_input_valid = io_input_valid; // @[port.scala 67:19]
  assign exponentArrayInHsk_io_input_bits_0_x_0 = io_input_bits_x_0; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_1 = io_input_bits_x_1; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_2 = io_input_bits_x_2; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_3 = io_input_bits_x_3; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_4 = io_input_bits_x_4; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_5 = io_input_bits_x_5; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_6 = io_input_bits_x_6; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_7 = io_input_bits_x_7; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_8 = io_input_bits_x_8; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_9 = io_input_bits_x_9; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_10 = io_input_bits_x_10; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_11 = io_input_bits_x_11; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_12 = io_input_bits_x_12; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_13 = io_input_bits_x_13; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_14 = io_input_bits_x_14; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_x_15 = io_input_bits_x_15; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_0_last = io_input_bits_last; // @[port.scala 65:27]
  assign exponentArrayInHsk_io_input_bits_1_x_0 = io_input_bits_x_0; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_1 = io_input_bits_x_1; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_2 = io_input_bits_x_2; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_3 = io_input_bits_x_3; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_4 = io_input_bits_x_4; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_5 = io_input_bits_x_5; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_6 = io_input_bits_x_6; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_7 = io_input_bits_x_7; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_8 = io_input_bits_x_8; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_9 = io_input_bits_x_9; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_10 = io_input_bits_x_10; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_11 = io_input_bits_x_11; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_12 = io_input_bits_x_12; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_13 = io_input_bits_x_13; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_14 = io_input_bits_x_14; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_x_15 = io_input_bits_x_15; // @[port.scala 62:19]
  assign exponentArrayInHsk_io_input_bits_1_last = io_input_bits_last; // @[port.scala 65:27]
  assign exponentArrayInHsk_io_output_0_ready = exponentArrayInMux_io_input_0_ready; // @[softmax.scala 51:41]
  assign exponentArrayInHsk_io_output_1_ready = queue_io_enq_ready; // @[softmax.scala 52:41]
  assign exponentArrayInMux_io_input_0_valid = exponentArrayInHsk_io_output_0_valid; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_0 = exponentArrayInHsk_io_output_0_bits_x_0; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_1 = exponentArrayInHsk_io_output_0_bits_x_1; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_2 = exponentArrayInHsk_io_output_0_bits_x_2; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_3 = exponentArrayInHsk_io_output_0_bits_x_3; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_4 = exponentArrayInHsk_io_output_0_bits_x_4; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_5 = exponentArrayInHsk_io_output_0_bits_x_5; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_6 = exponentArrayInHsk_io_output_0_bits_x_6; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_7 = exponentArrayInHsk_io_output_0_bits_x_7; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_8 = exponentArrayInHsk_io_output_0_bits_x_8; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_9 = exponentArrayInHsk_io_output_0_bits_x_9; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_10 = exponentArrayInHsk_io_output_0_bits_x_10; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_11 = exponentArrayInHsk_io_output_0_bits_x_11; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_12 = exponentArrayInHsk_io_output_0_bits_x_12; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_13 = exponentArrayInHsk_io_output_0_bits_x_13; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_14 = exponentArrayInHsk_io_output_0_bits_x_14; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_x_15 = exponentArrayInHsk_io_output_0_bits_x_15; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_0_bits_last = exponentArrayInHsk_io_output_0_bits_last; // @[softmax.scala 51:41]
  assign exponentArrayInMux_io_input_1_valid = adder_io_output_valid; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_0 = adder_io_output_bits_x_0; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_1 = adder_io_output_bits_x_1; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_2 = adder_io_output_bits_x_2; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_3 = adder_io_output_bits_x_3; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_4 = adder_io_output_bits_x_4; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_5 = adder_io_output_bits_x_5; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_6 = adder_io_output_bits_x_6; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_7 = adder_io_output_bits_x_7; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_8 = adder_io_output_bits_x_8; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_9 = adder_io_output_bits_x_9; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_10 = adder_io_output_bits_x_10; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_11 = adder_io_output_bits_x_11; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_12 = adder_io_output_bits_x_12; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_13 = adder_io_output_bits_x_13; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_14 = adder_io_output_bits_x_14; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_x_15 = adder_io_output_bits_x_15; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_input_1_bits_last = adder_io_output_bits_last; // @[softmax.scala 53:25]
  assign exponentArrayInMux_io_sel = inPathSel; // @[softmax.scala 69:35]
  assign exponentArrayInMux_io_output_ready = exponentArray_io_input_ready; // @[softmax.scala 54:38]
  assign exponentArrayOutMux_io_input_valid = exponentArray_io_output_valid; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_0 = exponentArray_io_output_bits_x_0; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_1 = exponentArray_io_output_bits_x_1; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_2 = exponentArray_io_output_bits_x_2; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_3 = exponentArray_io_output_bits_x_3; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_4 = exponentArray_io_output_bits_x_4; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_5 = exponentArray_io_output_bits_x_5; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_6 = exponentArray_io_output_bits_x_6; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_7 = exponentArray_io_output_bits_x_7; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_8 = exponentArray_io_output_bits_x_8; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_9 = exponentArray_io_output_bits_x_9; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_10 = exponentArray_io_output_bits_x_10; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_11 = exponentArray_io_output_bits_x_11; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_12 = exponentArray_io_output_bits_x_12; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_13 = exponentArray_io_output_bits_x_13; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_14 = exponentArray_io_output_bits_x_14; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_x_15 = exponentArray_io_output_bits_x_15; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_input_bits_last = exponentArray_io_output_bits_last; // @[softmax.scala 57:33]
  assign exponentArrayOutMux_io_sel = outPathSel; // @[softmax.scala 71:36]
  assign exponentArrayOutMux_io_output_0_ready = adderTree_io_input_ready; // @[softmax.scala 58:42]
  assign exponentArrayOutMux_io_output_1_ready = io_output_ready; // @[softmax.scala 59:42]
  assign queue_clock = clock;
  assign queue_reset = rst;
  assign queue_io_enq_valid = exponentArrayInHsk_io_output_1_valid; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_0 = exponentArrayInHsk_io_output_1_bits_x_0; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_1 = exponentArrayInHsk_io_output_1_bits_x_1; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_2 = exponentArrayInHsk_io_output_1_bits_x_2; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_3 = exponentArrayInHsk_io_output_1_bits_x_3; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_4 = exponentArrayInHsk_io_output_1_bits_x_4; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_5 = exponentArrayInHsk_io_output_1_bits_x_5; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_6 = exponentArrayInHsk_io_output_1_bits_x_6; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_7 = exponentArrayInHsk_io_output_1_bits_x_7; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_8 = exponentArrayInHsk_io_output_1_bits_x_8; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_9 = exponentArrayInHsk_io_output_1_bits_x_9; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_10 = exponentArrayInHsk_io_output_1_bits_x_10; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_11 = exponentArrayInHsk_io_output_1_bits_x_11; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_12 = exponentArrayInHsk_io_output_1_bits_x_12; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_13 = exponentArrayInHsk_io_output_1_bits_x_13; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_14 = exponentArrayInHsk_io_output_1_bits_x_14; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_x_15 = exponentArrayInHsk_io_output_1_bits_x_15; // @[softmax.scala 52:41]
  assign queue_io_enq_bits_last = exponentArrayInHsk_io_output_1_bits_last; // @[softmax.scala 52:41]
  assign queue_io_deq_ready = queueOutHsk_io_input_0_ready; // @[softmax.scala 64:22]
  assign adder_clock = clock;
  assign adder_reset = rst;
  assign adder_io_input_valid = queueOutHsk_io_output_valid; // @[port.scala 24:19]
  assign adder_io_input_bits_x_0 = queueOutHsk_io_output_bits_0_x_0; // @[port.scala 20:37]
  assign adder_io_input_bits_x_1 = queueOutHsk_io_output_bits_0_x_1; // @[port.scala 20:37]
  assign adder_io_input_bits_x_2 = queueOutHsk_io_output_bits_0_x_2; // @[port.scala 20:37]
  assign adder_io_input_bits_x_3 = queueOutHsk_io_output_bits_0_x_3; // @[port.scala 20:37]
  assign adder_io_input_bits_x_4 = queueOutHsk_io_output_bits_0_x_4; // @[port.scala 20:37]
  assign adder_io_input_bits_x_5 = queueOutHsk_io_output_bits_0_x_5; // @[port.scala 20:37]
  assign adder_io_input_bits_x_6 = queueOutHsk_io_output_bits_0_x_6; // @[port.scala 20:37]
  assign adder_io_input_bits_x_7 = queueOutHsk_io_output_bits_0_x_7; // @[port.scala 20:37]
  assign adder_io_input_bits_x_8 = queueOutHsk_io_output_bits_0_x_8; // @[port.scala 20:37]
  assign adder_io_input_bits_x_9 = queueOutHsk_io_output_bits_0_x_9; // @[port.scala 20:37]
  assign adder_io_input_bits_x_10 = queueOutHsk_io_output_bits_0_x_10; // @[port.scala 20:37]
  assign adder_io_input_bits_x_11 = queueOutHsk_io_output_bits_0_x_11; // @[port.scala 20:37]
  assign adder_io_input_bits_x_12 = queueOutHsk_io_output_bits_0_x_12; // @[port.scala 20:37]
  assign adder_io_input_bits_x_13 = queueOutHsk_io_output_bits_0_x_13; // @[port.scala 20:37]
  assign adder_io_input_bits_x_14 = queueOutHsk_io_output_bits_0_x_14; // @[port.scala 20:37]
  assign adder_io_input_bits_x_15 = queueOutHsk_io_output_bits_0_x_15; // @[port.scala 20:37]
  assign adder_io_input_bits_x_16 = queueOutHsk_io_output_bits_1_x_0; // @[port.scala 20:37]
  assign adder_io_input_bits_x_17 = queueOutHsk_io_output_bits_1_x_1; // @[port.scala 20:37]
  assign adder_io_input_bits_x_18 = queueOutHsk_io_output_bits_1_x_2; // @[port.scala 20:37]
  assign adder_io_input_bits_x_19 = queueOutHsk_io_output_bits_1_x_3; // @[port.scala 20:37]
  assign adder_io_input_bits_x_20 = queueOutHsk_io_output_bits_1_x_4; // @[port.scala 20:37]
  assign adder_io_input_bits_x_21 = queueOutHsk_io_output_bits_1_x_5; // @[port.scala 20:37]
  assign adder_io_input_bits_x_22 = queueOutHsk_io_output_bits_1_x_6; // @[port.scala 20:37]
  assign adder_io_input_bits_x_23 = queueOutHsk_io_output_bits_1_x_7; // @[port.scala 20:37]
  assign adder_io_input_bits_x_24 = queueOutHsk_io_output_bits_1_x_8; // @[port.scala 20:37]
  assign adder_io_input_bits_x_25 = queueOutHsk_io_output_bits_1_x_9; // @[port.scala 20:37]
  assign adder_io_input_bits_x_26 = queueOutHsk_io_output_bits_1_x_10; // @[port.scala 20:37]
  assign adder_io_input_bits_x_27 = queueOutHsk_io_output_bits_1_x_11; // @[port.scala 20:37]
  assign adder_io_input_bits_x_28 = queueOutHsk_io_output_bits_1_x_12; // @[port.scala 20:37]
  assign adder_io_input_bits_x_29 = queueOutHsk_io_output_bits_1_x_13; // @[port.scala 20:37]
  assign adder_io_input_bits_x_30 = queueOutHsk_io_output_bits_1_x_14; // @[port.scala 20:37]
  assign adder_io_input_bits_x_31 = queueOutHsk_io_output_bits_1_x_15; // @[port.scala 20:37]
  assign adder_io_input_bits_last = queueOutHsk_io_output_bits_0_last; // @[port.scala 23:23]
  assign adder_io_output_ready = exponentArrayInMux_io_input_1_ready; // @[softmax.scala 53:25]
  assign adderTree_clock = clock;
  assign adderTree_reset = rst;
  assign adderTree_io_input_valid = exponentArrayOutMux_io_output_0_valid; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_0 = {{4{exponentArrayOutMux_io_output_0_bits_x_0[7]}},
    exponentArrayOutMux_io_output_0_bits_x_0}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_1 = {{4{exponentArrayOutMux_io_output_0_bits_x_1[7]}},
    exponentArrayOutMux_io_output_0_bits_x_1}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_2 = {{4{exponentArrayOutMux_io_output_0_bits_x_2[7]}},
    exponentArrayOutMux_io_output_0_bits_x_2}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_3 = {{4{exponentArrayOutMux_io_output_0_bits_x_3[7]}},
    exponentArrayOutMux_io_output_0_bits_x_3}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_4 = {{4{exponentArrayOutMux_io_output_0_bits_x_4[7]}},
    exponentArrayOutMux_io_output_0_bits_x_4}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_5 = {{4{exponentArrayOutMux_io_output_0_bits_x_5[7]}},
    exponentArrayOutMux_io_output_0_bits_x_5}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_6 = {{4{exponentArrayOutMux_io_output_0_bits_x_6[7]}},
    exponentArrayOutMux_io_output_0_bits_x_6}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_7 = {{4{exponentArrayOutMux_io_output_0_bits_x_7[7]}},
    exponentArrayOutMux_io_output_0_bits_x_7}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_8 = {{4{exponentArrayOutMux_io_output_0_bits_x_8[7]}},
    exponentArrayOutMux_io_output_0_bits_x_8}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_9 = {{4{exponentArrayOutMux_io_output_0_bits_x_9[7]}},
    exponentArrayOutMux_io_output_0_bits_x_9}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_10 = {{4{exponentArrayOutMux_io_output_0_bits_x_10[7]}},
    exponentArrayOutMux_io_output_0_bits_x_10}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_11 = {{4{exponentArrayOutMux_io_output_0_bits_x_11[7]}},
    exponentArrayOutMux_io_output_0_bits_x_11}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_12 = {{4{exponentArrayOutMux_io_output_0_bits_x_12[7]}},
    exponentArrayOutMux_io_output_0_bits_x_12}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_13 = {{4{exponentArrayOutMux_io_output_0_bits_x_13[7]}},
    exponentArrayOutMux_io_output_0_bits_x_13}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_14 = {{4{exponentArrayOutMux_io_output_0_bits_x_14[7]}},
    exponentArrayOutMux_io_output_0_bits_x_14}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_x_15 = {{4{exponentArrayOutMux_io_output_0_bits_x_15[7]}},
    exponentArrayOutMux_io_output_0_bits_x_15}; // @[softmax.scala 58:42]
  assign adderTree_io_input_bits_last = exponentArrayOutMux_io_output_0_bits_last; // @[softmax.scala 58:42]
  assign accumulator_clock = clock;
  assign accumulator_reset = rst;
  assign accumulator_io_input_valid = adderTree_io_output_valid; // @[softmax.scala 62:29]
  assign accumulator_io_input_bits_x_0 = adderTree_io_output_bits_x_0; // @[softmax.scala 62:29]
  assign accumulator_io_input_bits_last = adderTree_io_output_bits_last; // @[softmax.scala 62:29]
  assign logarithm_clock = clock;
  assign logarithm_reset = rst;
  assign logarithm_io_input_valid = accumulator_io_output_valid; // @[softmax.scala 63:31]
  assign logarithm_io_input_bits_x_0 = accumulator_io_output_bits_x_0; // @[softmax.scala 63:31]
  assign logarithm_io_input_bits_last = accumulator_io_output_bits_last; // @[softmax.scala 63:31]
  assign logarithm_io_output_ready = queueOutHsk_io_input_1_ready; // @[port.scala 46:19]
  assign queueOutHsk_io_input_0_valid = queue_io_deq_valid; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_0 = queue_io_deq_bits_x_0; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_1 = queue_io_deq_bits_x_1; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_2 = queue_io_deq_bits_x_2; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_3 = queue_io_deq_bits_x_3; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_4 = queue_io_deq_bits_x_4; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_5 = queue_io_deq_bits_x_5; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_6 = queue_io_deq_bits_x_6; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_7 = queue_io_deq_bits_x_7; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_8 = queue_io_deq_bits_x_8; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_9 = queue_io_deq_bits_x_9; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_10 = queue_io_deq_bits_x_10; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_11 = queue_io_deq_bits_x_11; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_12 = queue_io_deq_bits_x_12; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_13 = queue_io_deq_bits_x_13; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_14 = queue_io_deq_bits_x_14; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_x_15 = queue_io_deq_bits_x_15; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_0_bits_last = queue_io_deq_bits_last; // @[softmax.scala 64:22]
  assign queueOutHsk_io_input_1_valid = logarithm_io_output_valid; // @[port.scala 45:19]
  assign queueOutHsk_io_input_1_bits_x_0 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_1 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_2 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_3 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_4 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_5 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_6 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_7 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_8 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_9 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_10 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_11 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_12 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_13 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_14 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_input_1_bits_x_15 = logarithm_io_output_bits_x_0; // @[port.scala 41:15]
  assign queueOutHsk_io_output_ready = adder_io_input_ready; // @[port.scala 25:19]
  always @(posedge clock or posedge rst) begin
    if (rst) begin // @[Reg.scala 29:18]
      inPathSel <= 1'h0; // @[Reg.scala 29:22]
    end else if (inPathSelEn) begin // @[Reg.scala 28:20]
      inPathSel <= inPathSelNxt;
    end
  end
  always @(posedge clock or posedge rst) begin
    if (rst) begin // @[Reg.scala 29:18]
      outPathSel <= 1'h0; // @[Reg.scala 29:22]
    end else if (outPathSelEn) begin // @[Reg.scala 28:20]
      outPathSel <= outPathSelNxt;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inPathSel = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  outPathSel = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  if (rst) begin
    inPathSel = 1'h0;
  end
  if (rst) begin
    outPathSel = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
